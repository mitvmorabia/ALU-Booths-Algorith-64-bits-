
module multiplier ( result, valid, opera1, opera2, muordi, clock, reset, start
 );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input muordi, clock, reset, start;
  output valid;
  wire   opera2_63, N34, n52, n53, n55, n56, n102, n104, n106, n108, n110,
         n112, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n991, n993, n994, n995, n997,
         n998, n1007, n1368, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1787, n1790, n1791, n1792, n1793, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1857, n1858, n1860, n1861, n1862,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2084, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2710, n2711, n2712, n2713, n2724, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784;
  wire   [63:0] res_not_wire;
  wire   [2:0] nst;
  wire   [31:0] i;
  tri   c_inop1;
  tri   c_inop2;
  tri   c_inres;
  assign opera2_63 = opera2[63];

  CTSX2 A5 ( .A(1'b1), .E(n1007), .Z(c_inres) );
  CTSX2 A4 ( .A(1'b0), .E(n1787), .Z(c_inop2) );
  CTSX2 A3 ( .A(1'b1), .E(n2704), .Z(c_inop2) );
  CTSX2 A1 ( .A(1'b1), .E(n2777), .Z(c_inop1) );
  CIVX2 U1559 ( .A(c_inop2), .Z(n2452) );
  CAN3X2 U1594 ( .A(n53), .B(n1936), .C(n56), .Z(n1988) );
  CAN3X2 U1605 ( .A(i[11]), .B(n2023), .C(i[12]), .Z(n2028) );
  CAN3X2 U1606 ( .A(i[10]), .B(n2018), .C(i[9]), .Z(n2023) );
  CAN3X2 U1607 ( .A(i[7]), .B(n2013), .C(i[8]), .Z(n2018) );
  CAN3X2 U1608 ( .A(i[5]), .B(n2002), .C(i[6]), .Z(n2013) );
  CAN3X2 U1609 ( .A(i[3]), .B(n1999), .C(i[4]), .Z(n2002) );
  CIVX2 U1626 ( .A(n2445), .Z(n1734) );
  CIVX2 U1627 ( .A(n2358), .Z(n1735) );
  CIVX2 U1628 ( .A(n2443), .Z(n1736) );
  CIVX2 U1630 ( .A(n2441), .Z(n1738) );
  CIVX2 U1631 ( .A(n2439), .Z(n1739) );
  CIVX2 U1632 ( .A(n2437), .Z(n1740) );
  CIVX2 U1633 ( .A(n2363), .Z(n1741) );
  CIVX2 U1634 ( .A(n2435), .Z(n1742) );
  CIVX2 U1636 ( .A(n2433), .Z(n1744) );
  CIVX2 U1637 ( .A(n2431), .Z(n1745) );
  CIVX2 U1638 ( .A(n2429), .Z(n1746) );
  CIVX2 U1639 ( .A(n2368), .Z(n1747) );
  CIVX2 U1640 ( .A(n2427), .Z(n1748) );
  CIVX2 U1642 ( .A(n2425), .Z(n1750) );
  CIVX2 U1643 ( .A(n2423), .Z(n1751) );
  CIVX2 U1644 ( .A(n2421), .Z(n1752) );
  CIVX2 U1645 ( .A(n2373), .Z(n1753) );
  CIVX2 U1646 ( .A(n2419), .Z(n1754) );
  CIVX2 U1648 ( .A(n2417), .Z(n1756) );
  CIVX2 U1649 ( .A(n2415), .Z(n1757) );
  CIVX2 U1650 ( .A(n2413), .Z(n1758) );
  CIVX2 U1651 ( .A(n2378), .Z(n1759) );
  CIVX2 U1654 ( .A(n2409), .Z(n1762) );
  CIVX2 U1655 ( .A(n2407), .Z(n1763) );
  CIVX2 U1656 ( .A(n2405), .Z(n1764) );
  CIVX2 U1657 ( .A(n2403), .Z(n1765) );
  CIVX2 U1658 ( .A(n2401), .Z(n1766) );
  CIVX2 U1659 ( .A(n2399), .Z(n1767) );
  CIVX2 U1660 ( .A(n2397), .Z(n1768) );
  CIVX2 U1666 ( .A(n2603), .Z(n1774) );
  CIVX2 U1667 ( .A(n2591), .Z(n1775) );
  CIVX2 U1668 ( .A(n2579), .Z(n1776) );
  CIVX2 U1669 ( .A(n2567), .Z(n1777) );
  CIVX2 U1677 ( .A(n2495), .Z(n1783) );
  CIVX2 U1678 ( .A(n2483), .Z(n1784) );
  CIVX2 U1679 ( .A(n2471), .Z(n1785) );
  CIVX2 U1689 ( .A(n2082), .Z(n1795) );
  CIVX2 U1690 ( .A(n1992), .Z(n1796) );
  CIVX2 U1691 ( .A(n2705), .Z(n1797) );
  CIVX2 U1692 ( .A(reset), .Z(n1798) );
  CIVX2 U1693 ( .A(n1989), .Z(n1799) );
  CIVX2 U1694 ( .A(n2075), .Z(n1800) );
  CIVX2 U1695 ( .A(n2155), .Z(n1801) );
  CIVX2 U1696 ( .A(n1990), .Z(n1802) );
  CIVX2 U1697 ( .A(n53), .Z(n1803) );
  CIVX2 U1713 ( .A(nst[2]), .Z(n1819) );
  CIVX2 U1715 ( .A(result[30]), .Z(n1821) );
  CIVX2 U1716 ( .A(result[28]), .Z(n1822) );
  CIVX2 U1717 ( .A(result[26]), .Z(n1823) );
  CIVX2 U1718 ( .A(result[24]), .Z(n1824) );
  CIVX2 U1719 ( .A(result[22]), .Z(n1825) );
  CIVX2 U1720 ( .A(result[20]), .Z(n1826) );
  CIVX2 U1721 ( .A(result[18]), .Z(n1827) );
  CIVX2 U1722 ( .A(result[16]), .Z(n1828) );
  CIVX2 U1723 ( .A(result[14]), .Z(n1829) );
  CIVX2 U1724 ( .A(result[12]), .Z(n1830) );
  CIVX2 U1725 ( .A(result[10]), .Z(n1831) );
  CIVX2 U1726 ( .A(result[6]), .Z(n1832) );
  CIVX2 U1727 ( .A(result[4]), .Z(n1833) );
  CIVX2 U1728 ( .A(result[2]), .Z(n1834) );
  CIVX2 U1729 ( .A(result[8]), .Z(n1835) );
  CIVX2 U1730 ( .A(result[29]), .Z(n1836) );
  CIVX2 U1731 ( .A(result[7]), .Z(n1837) );
  CIVX2 U1732 ( .A(result[5]), .Z(n1838) );
  CIVX2 U1733 ( .A(result[3]), .Z(n1839) );
  CIVX2 U1734 ( .A(result[1]), .Z(n1840) );
  CIVX2 U1735 ( .A(result[27]), .Z(n1841) );
  CIVX2 U1736 ( .A(result[25]), .Z(n1842) );
  CIVX2 U1737 ( .A(result[23]), .Z(n1843) );
  CIVX2 U1738 ( .A(result[21]), .Z(n1844) );
  CIVX2 U1739 ( .A(result[19]), .Z(n1845) );
  CIVX2 U1740 ( .A(result[17]), .Z(n1846) );
  CIVX2 U1741 ( .A(result[15]), .Z(n1847) );
  CIVX2 U1742 ( .A(result[13]), .Z(n1848) );
  CIVX2 U1743 ( .A(result[11]), .Z(n1849) );
  CIVX2 U1744 ( .A(result[9]), .Z(n1850) );
  CIVX2 U1745 ( .A(result[63]), .Z(n1851) );
  CIVX2 U1746 ( .A(n104), .Z(n1852) );
  CIVX2 U1747 ( .A(n108), .Z(n1853) );
  CIVX2 U1748 ( .A(result[0]), .Z(n1854) );
  CIVX2 U1749 ( .A(n112), .Z(n1855) );
  CIVX2 U1751 ( .A(n998), .Z(n1857) );
  CIVX2 U1752 ( .A(n997), .Z(n1858) );
  CIVX2 U1754 ( .A(n995), .Z(n1860) );
  CIVX2 U1755 ( .A(n994), .Z(n1861) );
  CIVX2 U1756 ( .A(n993), .Z(n1862) );
  CIVX2 U1758 ( .A(n991), .Z(n1864) );
  CIVX2 U1759 ( .A(i[24]), .Z(n1865) );
  CIVX2 U1760 ( .A(n1995), .Z(n1866) );
  CIVX2 U1761 ( .A(n2066), .Z(n1867) );
  CIVX2 U1762 ( .A(n2065), .Z(n1868) );
  CIVX2 U1763 ( .A(n2056), .Z(n1869) );
  CIVX2 U1764 ( .A(n2163), .Z(n1870) );
  CIVX2 U1766 ( .A(i[27]), .Z(n1872) );
  CIVX2 U1767 ( .A(i[28]), .Z(n1873) );
  CIVX2 U1768 ( .A(i[20]), .Z(n1874) );
  CIVX2 U1769 ( .A(n2055), .Z(n1875) );
  CIVX2 U1770 ( .A(n2046), .Z(n1876) );
  CIVX2 U1771 ( .A(i[25]), .Z(n1877) );
  CIVX2 U1772 ( .A(i[23]), .Z(n1878) );
  CIVX2 U1773 ( .A(i[21]), .Z(n1879) );
  CIVX2 U1774 ( .A(i[31]), .Z(n1880) );
  CIVX2 U1775 ( .A(n989), .Z(n1881) );
  CIVX2 U1776 ( .A(n988), .Z(n1882) );
  CIVX2 U1777 ( .A(n2628), .Z(n1883) );
  CIVX2 U1778 ( .A(n2045), .Z(n1884) );
  CIVX2 U1779 ( .A(i[18]), .Z(n1885) );
  CIVX2 U1780 ( .A(i[17]), .Z(n1886) );
  CIVX2 U1781 ( .A(i[29]), .Z(n1887) );
  CIVX2 U1782 ( .A(n987), .Z(n1888) );
  CIVX2 U1783 ( .A(n2616), .Z(n1889) );
  CIVX2 U1786 ( .A(n986), .Z(n1892) );
  CIVX2 U1787 ( .A(i[19]), .Z(n1893) );
  CIVX2 U1788 ( .A(n2036), .Z(n1894) );
  CIVX2 U1789 ( .A(i[16]), .Z(n1895) );
  CIVX2 U1790 ( .A(n985), .Z(n1896) );
  CIVX2 U1791 ( .A(i[12]), .Z(n1897) );
  CIVX2 U1792 ( .A(n2035), .Z(n1898) );
  CIVX2 U1793 ( .A(i[15]), .Z(n1899) );
  CIVX2 U1794 ( .A(i[14]), .Z(n1900) );
  CIVX2 U1795 ( .A(i[13]), .Z(n1901) );
  CIVX2 U1796 ( .A(n984), .Z(n1902) );
  CIVX2 U1798 ( .A(n2568), .Z(n1904) );
  CIVX2 U1800 ( .A(n983), .Z(n1906) );
  CIVX2 U1801 ( .A(n2544), .Z(n1907) );
  CIVX2 U1802 ( .A(n982), .Z(n1908) );
  CIVX2 U1803 ( .A(n981), .Z(n1909) );
  CIVX2 U1805 ( .A(n2532), .Z(n1911) );
  CIVX2 U1806 ( .A(n2520), .Z(n1912) );
  CIVX2 U1807 ( .A(n2508), .Z(n1913) );
  CIVX2 U1808 ( .A(i[10]), .Z(n1914) );
  CIVX2 U1809 ( .A(i[8]), .Z(n1915) );
  CIVX2 U1810 ( .A(i[9]), .Z(n1916) );
  CIVX2 U1811 ( .A(i[7]), .Z(n1917) );
  CIVX2 U1812 ( .A(n979), .Z(n1918) );
  CIVX2 U1813 ( .A(n978), .Z(n1919) );
  CIVX2 U1814 ( .A(i[11]), .Z(n1920) );
  CIVX2 U1815 ( .A(n977), .Z(n1921) );
  CIVX2 U1816 ( .A(n2496), .Z(n1922) );
  CIVX2 U1817 ( .A(i[4]), .Z(n1923) );
  CIVX2 U1818 ( .A(i[6]), .Z(n1924) );
  CIVX2 U1819 ( .A(i[3]), .Z(n1925) );
  CIVX2 U1820 ( .A(i[5]), .Z(n1926) );
  CIVX2 U1824 ( .A(i[2]), .Z(n1930) );
  CIVX2 U1825 ( .A(n975), .Z(n1931) );
  CIVX2 U1826 ( .A(n2472), .Z(n1932) );
  CIVX2 U1827 ( .A(n974), .Z(n1933) );
  CIVX2 U1828 ( .A(n2460), .Z(n1934) );
  CIVX2 U1831 ( .A(res_not_wire[62]), .Z(n1937) );
  CIVX2 U1832 ( .A(res_not_wire[60]), .Z(n1938) );
  CIVX2 U1833 ( .A(res_not_wire[58]), .Z(n1939) );
  CIVX2 U1834 ( .A(res_not_wire[56]), .Z(n1940) );
  CIVX2 U1835 ( .A(res_not_wire[54]), .Z(n1941) );
  CIVX2 U1836 ( .A(res_not_wire[52]), .Z(n1942) );
  CIVX2 U1837 ( .A(res_not_wire[50]), .Z(n1943) );
  CIVX2 U1838 ( .A(res_not_wire[48]), .Z(n1944) );
  CIVX2 U1839 ( .A(res_not_wire[46]), .Z(n1945) );
  CIVX2 U1840 ( .A(res_not_wire[44]), .Z(n1946) );
  CIVX2 U1841 ( .A(res_not_wire[42]), .Z(n1947) );
  CIVX2 U1842 ( .A(res_not_wire[40]), .Z(n1948) );
  CIVX2 U1843 ( .A(res_not_wire[38]), .Z(n1949) );
  CIVX2 U1844 ( .A(res_not_wire[36]), .Z(n1950) );
  CIVX2 U1845 ( .A(res_not_wire[34]), .Z(n1951) );
  CIVX2 U1847 ( .A(res_not_wire[26]), .Z(n1953) );
  CIVX2 U1849 ( .A(res_not_wire[22]), .Z(n1955) );
  CIVX2 U1851 ( .A(res_not_wire[18]), .Z(n1957) );
  CIVX2 U1853 ( .A(res_not_wire[14]), .Z(n1959) );
  CIVX2 U1855 ( .A(res_not_wire[10]), .Z(n1961) );
  CIVX2 U1857 ( .A(res_not_wire[6]), .Z(n1963) );
  CIVX2 U1858 ( .A(n2701), .Z(n1964) );
  CIVX2 U1859 ( .A(res_not_wire[2]), .Z(n1965) );
  CIVX2 U1860 ( .A(res_not_wire[32]), .Z(n1966) );
  CIVX2 U1861 ( .A(res_not_wire[30]), .Z(n1967) );
  CIVX2 U1863 ( .A(result[60]), .Z(n1969) );
  CIVX2 U1864 ( .A(result[58]), .Z(n1970) );
  CIVX2 U1865 ( .A(result[56]), .Z(n1971) );
  CIVX2 U1866 ( .A(result[54]), .Z(n1972) );
  CIVX2 U1867 ( .A(result[52]), .Z(n1973) );
  CIVX2 U1868 ( .A(result[50]), .Z(n1974) );
  CIVX2 U1869 ( .A(result[48]), .Z(n1975) );
  CIVX2 U1870 ( .A(result[46]), .Z(n1976) );
  CIVX2 U1871 ( .A(result[44]), .Z(n1977) );
  CIVX2 U1872 ( .A(result[42]), .Z(n1978) );
  CIVX2 U1873 ( .A(result[40]), .Z(n1979) );
  CIVX2 U1874 ( .A(result[38]), .Z(n1980) );
  CIVX2 U1875 ( .A(result[36]), .Z(n1981) );
  CIVX2 U1876 ( .A(result[34]), .Z(n1982) );
  CIVX2 U1877 ( .A(result[62]), .Z(n1983) );
  CIVX2 U1878 ( .A(result[61]), .Z(n1984) );
  CIVX2 U1879 ( .A(i[0]), .Z(n1985) );
  CIVX2 U1880 ( .A(i[1]), .Z(n1986) );
  COAN1X1 U1881 ( .A(i[0]), .B(n2745), .C(n2744), .Z(n2003) );
  COAN1X1 U1882 ( .A(n1999), .B(n1994), .C(n2743), .Z(n1996) );
  COAN1X1 U1883 ( .A(n2002), .B(n2745), .C(n1993), .Z(n2000) );
  COAN1X1 U1884 ( .A(n2013), .B(n1994), .C(n2744), .Z(n2011) );
  COAN1X1 U1885 ( .A(n2018), .B(n2745), .C(n2743), .Z(n2016) );
  COAN1X1 U1886 ( .A(n2023), .B(n1994), .C(n1993), .Z(n2021) );
  COAN1X1 U1887 ( .A(n2028), .B(n2745), .C(n2744), .Z(n2026) );
  COR4X1 U1888 ( .A(n1899), .B(n2745), .C(i[16]), .D(n2035), .Z(n2034) );
  COAN1X1 U1889 ( .A(n1898), .B(n1994), .C(n2743), .Z(n2031) );
  COR4X1 U1890 ( .A(n1893), .B(n1994), .C(i[20]), .D(n2045), .Z(n2044) );
  COAN1X1 U1891 ( .A(n1884), .B(n2745), .C(n1993), .Z(n2041) );
  COR4X1 U1892 ( .A(n1994), .B(n1879), .C(n2046), .D(i[22]), .Z(n2050) );
  COR4X1 U1893 ( .A(n1878), .B(n2745), .C(i[24]), .D(n2055), .Z(n2054) );
  COAN1X1 U1894 ( .A(n1875), .B(n1994), .C(n1993), .Z(n2051) );
  COR4X1 U1895 ( .A(n2745), .B(n1877), .C(n2056), .D(i[26]), .Z(n2060) );
  COR4X1 U1896 ( .A(n1872), .B(n1994), .C(i[28]), .D(n2065), .Z(n2064) );
  COAN1X1 U1897 ( .A(n1868), .B(n1994), .C(n1993), .Z(n2061) );
  COR4X1 U1898 ( .A(n1994), .B(n1887), .C(n2066), .D(i[30]), .Z(n2070) );
  CAOR2X1 U1899 ( .A(n2769), .B(n1801), .C(valid), .D(n2657), .Z(n923) );
  CAOR1X1 U1900 ( .A(n2354), .B(n2353), .C(n1983), .Z(n2356) );
  CND2IX1 U1901 ( .B(n2153), .A(n2156), .Z(n2391) );
  COAN1X1 U1902 ( .A(n1769), .B(n2396), .C(n2397), .Z(n2387) );
  COAN1X1 U1903 ( .A(n1767), .B(n2400), .C(n2401), .Z(n2385) );
  COAN1X1 U1904 ( .A(n1765), .B(n2404), .C(n2405), .Z(n2383) );
  COAN1X1 U1905 ( .A(n1763), .B(n2408), .C(n2409), .Z(n2381) );
  COAN1X1 U1906 ( .A(n1757), .B(n2416), .C(n2417), .Z(n2376) );
  COAN1X1 U1907 ( .A(n1751), .B(n2424), .C(n2425), .Z(n2371) );
  COAN1X1 U1908 ( .A(n1745), .B(n2432), .C(n2433), .Z(n2366) );
  COAN1X1 U1909 ( .A(n1739), .B(n2440), .C(n2441), .Z(n2361) );
  CND2IX1 U1910 ( .B(n2627), .A(n2640), .Z(n2639) );
  COR8X1 U1911 ( .A(n2648), .B(n2649), .C(n2650), .D(n2646), .E(n2155), .F(
        i[1]), .G(i[0]), .H(n2651), .Z(n2075) );
  COR4X1 U1912 ( .A(n2650), .B(n2649), .C(n2648), .D(i[5]), .Z(n2652) );
  COR8X1 U1913 ( .A(i[13]), .B(i[12]), .C(i[10]), .D(n2653), .E(i[28]), .F(
        i[27]), .G(i[25]), .H(n2654), .Z(n2650) );
  COR8X1 U1914 ( .A(i[20]), .B(i[17]), .C(i[22]), .D(i[21]), .E(i[26]), .F(
        i[24]), .G(i[9]), .H(i[30]), .Z(n2649) );
  CAN4X1 U1915 ( .A(n56), .B(n53), .C(n1368), .D(reset), .Z(n2078) );
  COR2X1 U1916 ( .A(n2707), .B(n2708), .Z(n52) );
  CFD1QXL \nst_reg[2]  ( .D(n921), .CP(clock), .Q(nst[2]) );
  CFD1QXL \nst_reg[0]  ( .D(n2687), .CP(clock), .Q(nst[0]) );
  CFD1XL \res_not_reg[61]  ( .D(n858), .CP(clock), .QN(n104) );
  CFD1QXL \result_reg[63]  ( .D(n919), .CP(clock), .Q(result[63]) );
  CFD1QXL \res_not_reg[62]  ( .D(n857), .CP(clock), .Q(res_not_wire[62]) );
  CFD1XL \result_reg[31]  ( .D(n794), .CP(clock), .Q(result[31]), .QN(n2684)
         );
  CFD1XL \res_not_reg[63]  ( .D(n793), .CP(clock), .QN(n102) );
  CFD1QXL \result_reg[30]  ( .D(n795), .CP(clock), .Q(result[30]) );
  CFD1QXL \result_reg[28]  ( .D(n797), .CP(clock), .Q(result[28]) );
  CFD1QXL \result_reg[26]  ( .D(n799), .CP(clock), .Q(result[26]) );
  CFD1QXL \result_reg[24]  ( .D(n801), .CP(clock), .Q(result[24]) );
  CFD1QXL \result_reg[22]  ( .D(n803), .CP(clock), .Q(result[22]) );
  CFD1QXL \result_reg[20]  ( .D(n805), .CP(clock), .Q(result[20]) );
  CFD1QXL \result_reg[18]  ( .D(n807), .CP(clock), .Q(result[18]) );
  CFD1QXL \result_reg[16]  ( .D(n809), .CP(clock), .Q(result[16]) );
  CFD1QXL \result_reg[14]  ( .D(n811), .CP(clock), .Q(result[14]) );
  CFD1QXL \result_reg[12]  ( .D(n813), .CP(clock), .Q(result[12]) );
  CFD1QXL \result_reg[10]  ( .D(n815), .CP(clock), .Q(result[10]) );
  CFD1QXL \result_reg[6]  ( .D(n819), .CP(clock), .Q(result[6]) );
  CFD1QXL \result_reg[4]  ( .D(n821), .CP(clock), .Q(result[4]) );
  CFD1QXL \result_reg[2]  ( .D(n823), .CP(clock), .Q(result[2]) );
  CFD1QXL \result_reg[8]  ( .D(n817), .CP(clock), .Q(result[8]) );
  CFD1QXL \result_reg[29]  ( .D(n796), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[7]  ( .D(n818), .CP(clock), .Q(result[7]) );
  CFD1QXL \result_reg[5]  ( .D(n820), .CP(clock), .Q(result[5]) );
  CFD1QXL \result_reg[3]  ( .D(n822), .CP(clock), .Q(result[3]) );
  CFD1QXL \result_reg[1]  ( .D(n824), .CP(clock), .Q(result[1]) );
  CFD1QXL \result_reg[27]  ( .D(n798), .CP(clock), .Q(result[27]) );
  CFD1QXL \result_reg[25]  ( .D(n800), .CP(clock), .Q(result[25]) );
  CFD1QXL \result_reg[23]  ( .D(n802), .CP(clock), .Q(result[23]) );
  CFD1QXL \result_reg[21]  ( .D(n804), .CP(clock), .Q(result[21]) );
  CFD1QXL \result_reg[19]  ( .D(n806), .CP(clock), .Q(result[19]) );
  CFD1QXL \result_reg[17]  ( .D(n808), .CP(clock), .Q(result[17]) );
  CFD1QXL \result_reg[15]  ( .D(n810), .CP(clock), .Q(result[15]) );
  CFD1QXL \result_reg[13]  ( .D(n812), .CP(clock), .Q(result[13]) );
  CFD1QXL \result_reg[11]  ( .D(n814), .CP(clock), .Q(result[11]) );
  CFD1QXL \result_reg[9]  ( .D(n816), .CP(clock), .Q(result[9]) );
  CFD1QXL \res_not_reg[60]  ( .D(n859), .CP(clock), .Q(res_not_wire[60]) );
  CFD1XL \res_not_reg[57]  ( .D(n862), .CP(clock), .QN(n108) );
  CFD1XL \res_not_reg[53]  ( .D(n866), .CP(clock), .QN(n112) );
  CFD1QXL \res_not_reg[58]  ( .D(n861), .CP(clock), .Q(res_not_wire[58]) );
  CFD1QXL \res_not_reg[54]  ( .D(n865), .CP(clock), .Q(res_not_wire[54]) );
  CFD1QXL \res_not_reg[56]  ( .D(n863), .CP(clock), .Q(res_not_wire[56]) );
  CFD1QXL \res_not_reg[52]  ( .D(n867), .CP(clock), .Q(res_not_wire[52]) );
  CFD1XL \res_not_reg[59]  ( .D(n860), .CP(clock), .QN(n106) );
  CFD1XL \res_not_reg[55]  ( .D(n864), .CP(clock), .QN(n110) );
  CFD1QXL \result_reg[62]  ( .D(n826), .CP(clock), .Q(result[62]) );
  CFD1QXL \result_reg[0]  ( .D(n825), .CP(clock), .Q(result[0]) );
  CFD1QXL \result_reg[60]  ( .D(n828), .CP(clock), .Q(result[60]) );
  CFD1QXL \result_reg[61]  ( .D(n827), .CP(clock), .Q(result[61]) );
  CFD1XL \res_not_reg[47]  ( .D(n872), .CP(clock), .QN(n2679) );
  CFD1XL \res_not_reg[51]  ( .D(n868), .CP(clock), .Q(n998) );
  CFD1QXL \res_not_reg[50]  ( .D(n869), .CP(clock), .Q(res_not_wire[50]) );
  CFD1QXL \res_not_reg[46]  ( .D(n873), .CP(clock), .Q(res_not_wire[46]) );
  CFD1XL \res_not_reg[49]  ( .D(n870), .CP(clock), .Q(n997) );
  CFD1XL \res_not_reg[45]  ( .D(n874), .CP(clock), .Q(n995) );
  CFD1QXL \res_not_reg[48]  ( .D(n871), .CP(clock), .Q(res_not_wire[48]) );
  CFD1QXL \res_not_reg[44]  ( .D(n875), .CP(clock), .Q(res_not_wire[44]) );
  CFD1QXL \result_reg[56]  ( .D(n832), .CP(clock), .Q(result[56]) );
  CFD1XL \result_reg[59]  ( .D(n829), .CP(clock), .Q(result[59]), .QN(n2683)
         );
  CFD1XL \result_reg[57]  ( .D(n831), .CP(clock), .Q(result[57]), .QN(n2682)
         );
  CFD1QXL \result_reg[58]  ( .D(n830), .CP(clock), .Q(result[58]) );
  CFD1QXL \i_reg[31]  ( .D(n955), .CP(clock), .Q(i[31]) );
  CFD1XL \res_not_reg[43]  ( .D(n876), .CP(clock), .QN(n2676) );
  CFD1XL \res_not_reg[39]  ( .D(n880), .CP(clock), .QN(n2671) );
  CFD4QXL \cst_reg[1]  ( .D(n52), .CP(clock), .SD(n1798), .Q(n53) );
  CFD1QXL \i_reg[19]  ( .D(n935), .CP(clock), .Q(i[19]) );
  CFD1QXL \i_reg[16]  ( .D(n938), .CP(clock), .Q(i[16]) );
  CFD4QXL \cst_reg[0]  ( .D(n55), .CP(clock), .SD(n1798), .Q(n56) );
  CFD1QXL \res_not_reg[42]  ( .D(n877), .CP(clock), .Q(res_not_wire[42]) );
  CFD1QXL \res_not_reg[38]  ( .D(n881), .CP(clock), .Q(res_not_wire[38]) );
  CFD1XL \res_not_reg[41]  ( .D(n878), .CP(clock), .Q(n994) );
  CFD1XL \res_not_reg[37]  ( .D(n882), .CP(clock), .Q(n993) );
  CFD1QXL \res_not_reg[40]  ( .D(n879), .CP(clock), .Q(res_not_wire[40]) );
  CFD1QXL \res_not_reg[36]  ( .D(n883), .CP(clock), .Q(res_not_wire[36]) );
  CFD1QXL \result_reg[52]  ( .D(n836), .CP(clock), .Q(result[52]) );
  CFD1XL \result_reg[55]  ( .D(n833), .CP(clock), .Q(result[55]), .QN(n2681)
         );
  CFD1XL \result_reg[53]  ( .D(n835), .CP(clock), .Q(result[53]), .QN(n2678)
         );
  CFD1QXL \result_reg[54]  ( .D(n834), .CP(clock), .Q(result[54]) );
  CFD1XL \res_not_reg[35]  ( .D(n884), .CP(clock), .Q(n991) );
  CFD1XL \res_not_reg[33]  ( .D(n886), .CP(clock), .QN(n2667) );
  CFD1QXL \i_reg[10]  ( .D(n944), .CP(clock), .Q(i[10]) );
  CFD1QXL \i_reg[12]  ( .D(n942), .CP(clock), .Q(i[12]) );
  CFD1QXL \i_reg[23]  ( .D(n931), .CP(clock), .Q(i[23]) );
  CFD1QXL \i_reg[15]  ( .D(n939), .CP(clock), .Q(i[15]) );
  CFD1QXL \i_reg[14]  ( .D(n940), .CP(clock), .Q(i[14]) );
  CFD1QXL \i_reg[27]  ( .D(n927), .CP(clock), .Q(i[27]) );
  CFD1QXL \i_reg[11]  ( .D(n943), .CP(clock), .Q(i[11]) );
  CFD1QXL \i_reg[9]  ( .D(n945), .CP(clock), .Q(i[9]) );
  CFD1QXL \i_reg[20]  ( .D(n934), .CP(clock), .Q(i[20]) );
  CFD1QXL \i_reg[24]  ( .D(n930), .CP(clock), .Q(i[24]) );
  CFD1QXL \res_not_reg[32]  ( .D(n887), .CP(clock), .Q(res_not_wire[32]) );
  CFD1QXL \i_reg[28]  ( .D(n926), .CP(clock), .Q(i[28]) );
  CFD1QXL \res_not_reg[34]  ( .D(n885), .CP(clock), .Q(res_not_wire[34]) );
  CFD1QXL \i_reg[13]  ( .D(n941), .CP(clock), .Q(i[13]) );
  CFD1QXL \i_reg[29]  ( .D(n925), .CP(clock), .Q(i[29]) );
  CFD1QXL \i_reg[30]  ( .D(n924), .CP(clock), .Q(i[30]) );
  CFD1QXL \i_reg[22]  ( .D(n932), .CP(clock), .Q(i[22]) );
  CFD1QXL \i_reg[25]  ( .D(n929), .CP(clock), .Q(i[25]) );
  CFD1QXL \i_reg[26]  ( .D(n928), .CP(clock), .Q(i[26]) );
  CFD1QXL \i_reg[21]  ( .D(n933), .CP(clock), .Q(i[21]) );
  CFD1QXL \i_reg[18]  ( .D(n936), .CP(clock), .Q(i[18]) );
  CFD1QXL \i_reg[17]  ( .D(n937), .CP(clock), .Q(i[17]) );
  CFD1QXL \result_reg[48]  ( .D(n840), .CP(clock), .Q(result[48]) );
  CFD1XL \result_reg[51]  ( .D(n837), .CP(clock), .Q(result[51]), .QN(n2675)
         );
  CFD1XL \result_reg[49]  ( .D(n839), .CP(clock), .Q(result[49]), .QN(n2674)
         );
  CFD1QXL \result_reg[50]  ( .D(n838), .CP(clock), .Q(result[50]) );
  CFD1QXL \i_reg[8]  ( .D(n946), .CP(clock), .Q(i[8]) );
  CFD1QXL \i_reg[4]  ( .D(n949), .CP(clock), .Q(i[4]) );
  CFD1QXL \i_reg[6]  ( .D(n948), .CP(clock), .Q(i[6]) );
  CFD1QXL \i_reg[7]  ( .D(n947), .CP(clock), .Q(i[7]) );
  CFD1QXL \i_reg[3]  ( .D(n954), .CP(clock), .Q(i[3]) );
  CFD1QXL \i_reg[5]  ( .D(n953), .CP(clock), .Q(i[5]) );
  CFD1XL \res_not_reg[31]  ( .D(n888), .CP(clock), .Q(n989) );
  CFD1XL \result_reg[47]  ( .D(n841), .CP(clock), .Q(result[47]), .QN(n2670)
         );
  CFD1XL \result_reg[45]  ( .D(n843), .CP(clock), .Q(result[45]), .QN(n2665)
         );
  CFD1QXL \res_not_reg[30]  ( .D(n889), .CP(clock), .Q(res_not_wire[30]) );
  CFD1QXL \result_reg[46]  ( .D(n842), .CP(clock), .Q(result[46]) );
  CFD1QXL \i_reg[2]  ( .D(n950), .CP(clock), .Q(i[2]) );
  CFD1QXL \i_reg[1]  ( .D(n951), .CP(clock), .Q(i[1]) );
  CFD1QXL \i_reg[0]  ( .D(n952), .CP(clock), .Q(i[0]) );
  CFD1QXL \result_reg[42]  ( .D(n846), .CP(clock), .Q(result[42]) );
  CFD1QXL \result_reg[44]  ( .D(n844), .CP(clock), .Q(result[44]) );
  CFD1XL \result_reg[43]  ( .D(n845), .CP(clock), .Q(result[43]), .QN(n2666)
         );
  CFD1XL \result_reg[41]  ( .D(n847), .CP(clock), .Q(result[41]), .QN(n2662)
         );
  CFD1XL \result_reg[39]  ( .D(n849), .CP(clock), .Q(result[39]), .QN(n2663)
         );
  CFD1XL \result_reg[37]  ( .D(n851), .CP(clock), .Q(result[37]), .QN(n2661)
         );
  CFD1QXL \result_reg[38]  ( .D(n850), .CP(clock), .Q(result[38]) );
  CFD1QXL \result_reg[40]  ( .D(n848), .CP(clock), .Q(result[40]) );
  CFD1QXL \result_reg[32]  ( .D(n856), .CP(clock), .Q(result[32]) );
  CFD1QXL \res_not_reg[6]  ( .D(n913), .CP(clock), .Q(res_not_wire[6]) );
  CFD1QXL \result_reg[34]  ( .D(n854), .CP(clock), .Q(result[34]) );
  CFD1XL \result_reg[35]  ( .D(n853), .CP(clock), .Q(result[35]), .QN(n2660)
         );
  CFD1QXL \result_reg[36]  ( .D(n852), .CP(clock), .Q(result[36]) );
  CFD1XL \result_reg[33]  ( .D(n855), .CP(clock), .Q(result[33]), .QN(n2659)
         );
  CFD1XL \res_not_reg[7]  ( .D(n912), .CP(clock), .Q(n977) );
  CFD1XL \res_not_reg[3]  ( .D(n916), .CP(clock), .Q(n975) );
  CFD1QXL \res_not_reg[2]  ( .D(n917), .CP(clock), .Q(res_not_wire[2]) );
  CTSXL A2 ( .A(1'b0), .E(n2784), .Z(c_inop1) );
  CFD1X1 \res_not_reg[5]  ( .D(n914), .CP(clock), .Q(n976) );
  CFD1X1 \res_not_reg[1]  ( .D(n2702), .CP(clock), .Q(n974) );
  CFD1X1 sign_reg ( .D(n2703), .CP(clock), .Q(n1007), .QN(n1935) );
  CTSX1 A6 ( .A(1'b0), .E(n1935), .Z(c_inres) );
  CFD1QXL \res_not_reg[26]  ( .D(n893), .CP(clock), .Q(res_not_wire[26]) );
  CFD1QXL \res_not_reg[28]  ( .D(n891), .CP(clock), .Q(res_not_wire[28]) );
  CFD1XL \res_not_reg[29]  ( .D(n890), .CP(clock), .Q(n988) );
  CFD1XL \res_not_reg[27]  ( .D(n892), .CP(clock), .Q(n986) );
  CFD1QXL \res_not_reg[24]  ( .D(n895), .CP(clock), .Q(res_not_wire[24]) );
  CFD1QXL \res_not_reg[20]  ( .D(n899), .CP(clock), .Q(res_not_wire[20]) );
  CFD1QXL \res_not_reg[22]  ( .D(n897), .CP(clock), .Q(res_not_wire[22]) );
  CFD1QXL \res_not_reg[18]  ( .D(n901), .CP(clock), .Q(res_not_wire[18]) );
  CFD1XL \res_not_reg[23]  ( .D(n896), .CP(clock), .Q(n987) );
  CFD1XL \res_not_reg[25]  ( .D(n894), .CP(clock), .Q(n985) );
  CFD1XL \res_not_reg[19]  ( .D(n900), .CP(clock), .Q(n982) );
  CFD1XL \res_not_reg[21]  ( .D(n898), .CP(clock), .Q(n981) );
  CFD1QXL \res_not_reg[16]  ( .D(n903), .CP(clock), .Q(res_not_wire[16]) );
  CFD1QXL \res_not_reg[12]  ( .D(n907), .CP(clock), .Q(res_not_wire[12]) );
  CFD1QXL \res_not_reg[8]  ( .D(n911), .CP(clock), .Q(res_not_wire[8]) );
  CFD1QXL \res_not_reg[14]  ( .D(n905), .CP(clock), .Q(res_not_wire[14]) );
  CFD1QXL \res_not_reg[10]  ( .D(n909), .CP(clock), .Q(res_not_wire[10]) );
  CFD1XL \res_not_reg[17]  ( .D(n902), .CP(clock), .Q(n984) );
  CFD1XL \res_not_reg[15]  ( .D(n904), .CP(clock), .Q(n983) );
  CFD1XL \res_not_reg[11]  ( .D(n908), .CP(clock), .Q(n979) );
  CFD1XL \res_not_reg[13]  ( .D(n906), .CP(clock), .Q(n978) );
  CFD2XL \cst_reg[2]  ( .D(N34), .CP(clock), .CD(n1798), .Q(n1936), .QN(n1368)
         );
  CFD1QXL valid_reg ( .D(n923), .CP(clock), .Q(valid) );
  CFD1XL \nst_reg[1]  ( .D(n922), .CP(clock), .QN(n1820) );
  CFD1XL \res_not_reg[9]  ( .D(n2700), .CP(clock), .Q(n980), .QN(n2685) );
  CFD1QXL \res_not_reg[0]  ( .D(n920), .CP(clock), .Q(res_not_wire[0]) );
  CFD1QXL \res_not_reg[4]  ( .D(n915), .CP(clock), .Q(res_not_wire[4]) );
  CIVX1 U1917 ( .A(n2615), .Z(n1773) );
  CND3X1 U1918 ( .A(n993), .B(n2181), .C(res_not_wire[36]), .Z(n2196) );
  CNR3X2 U1919 ( .A(n1864), .B(n1870), .C(n1951), .Z(n2181) );
  CND3XL U1920 ( .A(n2283), .B(n1855), .C(res_not_wire[52]), .Z(n2297) );
  CND3XL U1921 ( .A(n2308), .B(n1853), .C(res_not_wire[56]), .Z(n2322) );
  CND3X1 U1922 ( .A(n979), .B(n1913), .C(res_not_wire[10]), .Z(n2520) );
  CND3X1 U1923 ( .A(n983), .B(n1911), .C(res_not_wire[14]), .Z(n2544) );
  CNR2X1 U1924 ( .A(n2472), .B(n2658), .Z(n2489) );
  CND3X1 U1925 ( .A(c_inres), .B(res_not_wire[0]), .C(n974), .Z(n2460) );
  CND3X1 U1926 ( .A(n980), .B(n1922), .C(res_not_wire[8]), .Z(n2508) );
  CND3X1 U1927 ( .A(n978), .B(n1912), .C(res_not_wire[12]), .Z(n2532) );
  CND3X1 U1928 ( .A(n984), .B(n1907), .C(res_not_wire[16]), .Z(n2556) );
  CND3X1 U1929 ( .A(n981), .B(n1904), .C(res_not_wire[20]), .Z(n2580) );
  CND3X1 U1930 ( .A(n985), .B(n1891), .C(res_not_wire[24]), .Z(n2604) );
  CND3X1 U1931 ( .A(n988), .B(n1889), .C(res_not_wire[28]), .Z(n2628) );
  CND3XL U1932 ( .A(n2333), .B(n1852), .C(res_not_wire[60]), .Z(n2086) );
  COND3XL U1933 ( .A(n2497), .B(n2747), .C(n2498), .D(n2499), .Z(n817) );
  COND3XL U1934 ( .A(n2473), .B(n2748), .C(n2474), .D(n2475), .Z(n821) );
  COND3XL U1935 ( .A(n2569), .B(n2746), .C(n2570), .D(n2571), .Z(n805) );
  COND3XL U1936 ( .A(n2593), .B(n2746), .C(n2594), .D(n2595), .Z(n801) );
  COND3XL U1937 ( .A(n2617), .B(n2746), .C(n2618), .D(n2619), .Z(n797) );
  CIVX2 U1938 ( .A(n2704), .Z(n1787) );
  CAN2X1 U1939 ( .A(n1988), .B(n2082), .Z(n2655) );
  COR3X2 U1940 ( .A(n2458), .B(n2453), .C(n2452), .Z(n2656) );
  CAN2X1 U1941 ( .A(n2645), .B(n2075), .Z(n2657) );
  COR2X1 U1942 ( .A(n1964), .B(n1928), .Z(n2658) );
  COR2X1 U1943 ( .A(n2513), .B(n2518), .Z(n2664) );
  COR2X1 U1944 ( .A(n1966), .B(n2667), .Z(n2668) );
  COR2X1 U1945 ( .A(n2525), .B(n2530), .Z(n2669) );
  COR2X1 U1946 ( .A(n1949), .B(n2671), .Z(n2672) );
  COR2X1 U1947 ( .A(n2549), .B(n2554), .Z(n2673) );
  COR2X1 U1948 ( .A(n1947), .B(n2676), .Z(n2677) );
  COR2X1 U1949 ( .A(n1945), .B(n2679), .Z(n2680) );
  CNIVXL U1950 ( .A(muordi), .Z(n2705) );
  CNIVX1 U1951 ( .A(n1797), .Z(n2686) );
  CNIVX1 U1952 ( .A(n957), .Z(n2687) );
  COND3X2 U1953 ( .A(n2082), .B(n2684), .C(n2634), .D(n2635), .Z(n794) );
  CEOXL U1954 ( .A(opera2[31]), .B(n2688), .Z(n2641) );
  CNIVX1 U1955 ( .A(opera2[30]), .Z(n2688) );
  CENX1 U1956 ( .A(opera2[29]), .B(n2704), .Z(n2626) );
  CNIVX1 U1957 ( .A(n2626), .Z(n2689) );
  CENX1 U1958 ( .A(opera2[7]), .B(n2704), .Z(n2494) );
  CNIVX1 U1959 ( .A(n2494), .Z(n2690) );
  CENX1 U1960 ( .A(opera2[5]), .B(n2704), .Z(n2482) );
  CNIVX1 U1961 ( .A(n2482), .Z(n2691) );
  CENX1 U1962 ( .A(opera2[3]), .B(n2704), .Z(n2470) );
  CNIVX1 U1963 ( .A(n2470), .Z(n2692) );
  CENXL U1964 ( .A(opera2[1]), .B(n2704), .Z(n2458) );
  CENX1 U1965 ( .A(opera2[27]), .B(n2704), .Z(n2614) );
  CNIVX1 U1966 ( .A(n2614), .Z(n2693) );
  CENX1 U1967 ( .A(opera2[25]), .B(n2704), .Z(n2602) );
  CNIVX1 U1968 ( .A(n2602), .Z(n2694) );
  CENX1 U1969 ( .A(opera2[23]), .B(n2704), .Z(n2590) );
  CNIVX1 U1970 ( .A(n2590), .Z(n2695) );
  CENX1 U1971 ( .A(opera2[21]), .B(n2704), .Z(n2578) );
  CNIVX1 U1972 ( .A(n2578), .Z(n2696) );
  CENX1 U1973 ( .A(opera2[19]), .B(n2704), .Z(n2566) );
  CNIVX1 U1974 ( .A(n2566), .Z(n2697) );
  CENXL U1975 ( .A(opera2[17]), .B(n2704), .Z(n2554) );
  CENX1 U1976 ( .A(opera2[15]), .B(n2704), .Z(n2542) );
  CNIVX1 U1977 ( .A(n2542), .Z(n2698) );
  CENXL U1978 ( .A(opera2[13]), .B(n2704), .Z(n2530) );
  CENXL U1979 ( .A(opera2[11]), .B(n2704), .Z(n2518) );
  CENX1 U1980 ( .A(opera2[9]), .B(n2704), .Z(n2506) );
  CNIVX1 U1981 ( .A(n2506), .Z(n2699) );
  COND1X1 U1982 ( .A(n106), .B(n2769), .C(n2145), .Z(n860) );
  COND1X1 U1983 ( .A(n110), .B(n2768), .C(n2141), .Z(n864) );
  COND3XL U1984 ( .A(n2353), .B(n2354), .C(n2355), .D(n2356), .Z(n2352) );
  CENXL U1985 ( .A(opera2[0]), .B(n2704), .Z(n2453) );
  CENXL U1986 ( .A(n2166), .B(n2167), .Z(n2165) );
  CNIVX1 U1987 ( .A(n910), .Z(n2700) );
  CIVXL U1988 ( .A(n976), .Z(n1928) );
  CNIVX1 U1989 ( .A(res_not_wire[4]), .Z(n2701) );
  CNIVX1 U1990 ( .A(n918), .Z(n2702) );
  CNIVX1 U1991 ( .A(n2706), .Z(n2703) );
  CNIVX4 U1992 ( .A(opera2_63), .Z(n2704) );
  CEOXL U1993 ( .A(n2704), .B(n2783), .Z(n1991) );
  CNIVX1 U1994 ( .A(n956), .Z(n2706) );
  COND2XL U1995 ( .A(n1796), .B(n1935), .C(n1991), .D(n1992), .Z(n956) );
  CDLY1XL U1996 ( .A(start), .Z(n2707) );
  CNR2XL U1997 ( .A(n2707), .B(n1819), .Z(N34) );
  CNIVX1 U1998 ( .A(n1820), .Z(n2708) );
  COR2X1 U1999 ( .A(n2664), .B(n1782), .Z(n1781) );
  CIVXL U2000 ( .A(n2507), .Z(n1782) );
  COR2X1 U2001 ( .A(n2669), .B(n1781), .Z(n1780) );
  COR2X1 U2002 ( .A(n2673), .B(n1779), .Z(n1778) );
  CIVXL U2003 ( .A(n2543), .Z(n1779) );
  CNR3XL U2004 ( .A(n2578), .B(n2573), .C(n1777), .Z(n2579) );
  CNR3XL U2005 ( .A(n2554), .B(n2549), .C(n1779), .Z(n2555) );
  CNR3XL U2006 ( .A(n2542), .B(n2537), .C(n1780), .Z(n2543) );
  CNR3XL U2007 ( .A(n2530), .B(n2525), .C(n1781), .Z(n2531) );
  CNR3XL U2008 ( .A(n2518), .B(n2513), .C(n1782), .Z(n2519) );
  CNR3XL U2009 ( .A(n2458), .B(n2453), .C(n2452), .Z(n2459) );
  CAN3X2 U2010 ( .A(n1772), .B(n1929), .C(n1792), .Z(n2710) );
  CNR2X1 U2011 ( .A(n2710), .B(n2636), .Z(n2635) );
  COND2XL U2012 ( .A(n2750), .B(n2637), .C(n2638), .D(n2639), .Z(n2636) );
  CNR3XL U2013 ( .A(n2566), .B(n2561), .C(n1778), .Z(n2567) );
  CENX1 U2014 ( .A(n2633), .B(n2627), .Z(n2632) );
  CNR2X1 U2015 ( .A(n2157), .B(n2668), .Z(n2163) );
  COND2X1 U2016 ( .A(n2663), .B(n2384), .C(n2201), .D(n2202), .Z(n2208) );
  COND2X1 U2017 ( .A(n2661), .B(n2386), .C(n2188), .D(n2189), .Z(n2194) );
  COND2X1 U2018 ( .A(n2683), .B(n2360), .C(n2327), .D(n2328), .Z(n2335) );
  COND2X1 U2019 ( .A(n1984), .B(n2357), .C(n1735), .D(n2340), .Z(n2347) );
  COND2X1 U2020 ( .A(n2665), .B(n2377), .C(n1759), .D(n2240), .Z(n2246) );
  COND2X1 U2021 ( .A(n2674), .B(n2372), .C(n1753), .D(n2265), .Z(n2271) );
  COND2X1 U2022 ( .A(n2678), .B(n2367), .C(n1747), .D(n2290), .Z(n2296) );
  COND2X1 U2023 ( .A(n2682), .B(n2362), .C(n1741), .D(n2315), .Z(n2321) );
  CNR2X1 U2024 ( .A(n2393), .B(n2392), .Z(n2166) );
  CAN2X1 U2025 ( .A(n2712), .B(n2713), .Z(n2156) );
  COND2X1 U2026 ( .A(n1971), .B(n2364), .C(n1743), .D(n2309), .Z(n2363) );
  COND2X1 U2027 ( .A(n1977), .B(n2379), .C(n1761), .D(n2234), .Z(n2378) );
  COND2X1 U2028 ( .A(n1975), .B(n2374), .C(n1755), .D(n2259), .Z(n2373) );
  COND2X1 U2029 ( .A(n1969), .B(n2359), .C(n1737), .D(n2334), .Z(n2358) );
  COND2X1 U2030 ( .A(n1973), .B(n2369), .C(n1749), .D(n2284), .Z(n2368) );
  CNR3XL U2031 ( .A(n2494), .B(n2488), .C(n1784), .Z(n2495) );
  CNR3XL U2032 ( .A(n2506), .B(n2501), .C(n1783), .Z(n2507) );
  CNR3XL U2033 ( .A(n2590), .B(n2585), .C(n1776), .Z(n2591) );
  CNR3XL U2034 ( .A(n2614), .B(n2609), .C(n1774), .Z(n2615) );
  CND3XL U2035 ( .A(n994), .B(n2207), .C(res_not_wire[40]), .Z(n2222) );
  CND3XL U2036 ( .A(n995), .B(n2233), .C(res_not_wire[44]), .Z(n2247) );
  CND3XL U2037 ( .A(n997), .B(n2258), .C(res_not_wire[48]), .Z(n2272) );
  CNR2X1 U2038 ( .A(n2247), .B(n2680), .Z(n2258) );
  CND2XL U2039 ( .A(n2392), .B(n2393), .Z(n2712) );
  CIVX2 U2040 ( .A(opera1[31]), .Z(n2784) );
  CIVXL U2041 ( .A(n2784), .Z(n2711) );
  CIVX2 U2042 ( .A(n2783), .Z(n2777) );
  CIVXL U2043 ( .A(n2166), .Z(n2713) );
  CIVX2 U2044 ( .A(n2156), .Z(n1770) );
  COND2X1 U2045 ( .A(n2662), .B(n2382), .C(n2214), .D(n2215), .Z(n2221) );
  CND2X1 U2046 ( .A(n1765), .B(n2404), .Z(n2405) );
  CND2X1 U2047 ( .A(n1767), .B(n2400), .Z(n2401) );
  CND2X1 U2048 ( .A(n1763), .B(n2408), .Z(n2409) );
  CND2X1 U2049 ( .A(n1769), .B(n2396), .Z(n2397) );
  CND2X1 U2050 ( .A(n1764), .B(n2406), .Z(n2407) );
  CND2X1 U2051 ( .A(n1766), .B(n2402), .Z(n2403) );
  CND2X1 U2052 ( .A(n1768), .B(n2398), .Z(n2399) );
  CNR3XL U2053 ( .A(n2626), .B(n2621), .C(n1773), .Z(n2627) );
  CNR3XL U2054 ( .A(n2482), .B(n2477), .C(n1785), .Z(n2483) );
  CNR3XL U2055 ( .A(n2470), .B(n2465), .C(n2656), .Z(n2471) );
  CNR3XL U2056 ( .A(n2602), .B(n2597), .C(n1775), .Z(n2603) );
  CNR2X1 U2057 ( .A(n2196), .B(n2672), .Z(n2207) );
  CND3X2 U2058 ( .A(n989), .B(n1883), .C(res_not_wire[30]), .Z(n2157) );
  CND3X2 U2059 ( .A(n975), .B(n1934), .C(res_not_wire[2]), .Z(n2472) );
  CENX1 U2060 ( .A(opera1[1]), .B(n2782), .Z(n2392) );
  CANR5CXL U2061 ( .A(result[34]), .B(n2389), .C(n2390), .Z(n2175) );
  CND2X1 U2062 ( .A(c_inop1), .B(n2644), .Z(n2393) );
  CIVX2 U2063 ( .A(opera1[31]), .Z(n2783) );
  CENX1 U2064 ( .A(n2208), .B(n2209), .Z(n2203) );
  CIVX1 U2065 ( .A(n2395), .Z(n1769) );
  CIVXL U2066 ( .A(n2411), .Z(n1760) );
  CEOXL U2067 ( .A(n2220), .B(n2221), .Z(n2219) );
  CANR4CXL U2068 ( .A(n2621), .B(n1773), .C(n2689), .D(n2627), .Z(n2625) );
  CEOXL U2069 ( .A(n1773), .B(n2621), .Z(n2620) );
  CANR4CXL U2070 ( .A(n2609), .B(n1774), .C(n2693), .D(n2615), .Z(n2613) );
  CANR4CXL U2071 ( .A(n2597), .B(n1775), .C(n2694), .D(n2603), .Z(n2601) );
  CEOXL U2072 ( .A(n2609), .B(n1774), .Z(n2608) );
  CANR4CXL U2073 ( .A(n2585), .B(n1776), .C(n2695), .D(n2591), .Z(n2589) );
  CEOXL U2074 ( .A(n1775), .B(n2597), .Z(n2596) );
  CIVX1 U2075 ( .A(n2235), .Z(n1761) );
  CIVX1 U2076 ( .A(n2260), .Z(n1755) );
  CIVX1 U2077 ( .A(n2310), .Z(n1743) );
  CIVX1 U2078 ( .A(n2335), .Z(n1737) );
  CIVX1 U2079 ( .A(n2285), .Z(n1749) );
  CANR4CXL U2080 ( .A(n2573), .B(n1777), .C(n2696), .D(n2579), .Z(n2577) );
  CANR4CXL U2081 ( .A(n2561), .B(n1778), .C(n2697), .D(n2567), .Z(n2565) );
  COND4CXL U2082 ( .A(n2166), .B(n2167), .C(n2394), .D(n2395), .Z(n2388) );
  CEOXL U2083 ( .A(n2585), .B(n1776), .Z(n2584) );
  CEOXL U2084 ( .A(n1777), .B(n2573), .Z(n2572) );
  CEOXL U2085 ( .A(n1735), .B(n2340), .Z(n2339) );
  CEOXL U2086 ( .A(n1741), .B(n2315), .Z(n2314) );
  CEOXL U2087 ( .A(n2327), .B(n2328), .Z(n2326) );
  CIVX1 U2088 ( .A(n2170), .Z(n1772) );
  CANR4CXL U2089 ( .A(n2549), .B(n1779), .C(n2554), .D(n2555), .Z(n2553) );
  CEOXL U2090 ( .A(n2561), .B(n1778), .Z(n2560) );
  CEOXL U2091 ( .A(n2302), .B(n2303), .Z(n2301) );
  CANR4CXL U2092 ( .A(n1772), .B(n2643), .C(n2344), .D(n1929), .Z(n2642) );
  CANR4CXL U2093 ( .A(n2537), .B(n1780), .C(n2698), .D(n2543), .Z(n2541) );
  CEOXL U2094 ( .A(n1779), .B(n2549), .Z(n2548) );
  CEOXL U2095 ( .A(n2277), .B(n2278), .Z(n2276) );
  CEOXL U2096 ( .A(n1747), .B(n2290), .Z(n2289) );
  CANR4CXL U2097 ( .A(n2525), .B(n1781), .C(n2530), .D(n2531), .Z(n2529) );
  CEOXL U2098 ( .A(n2537), .B(n1780), .Z(n2536) );
  CEOXL U2099 ( .A(n1753), .B(n2265), .Z(n2264) );
  CANR4CXL U2100 ( .A(n2513), .B(n1782), .C(n2518), .D(n2519), .Z(n2517) );
  CEOXL U2101 ( .A(n1781), .B(n2525), .Z(n2524) );
  CEOXL U2102 ( .A(n1759), .B(n2240), .Z(n2239) );
  CEOXL U2103 ( .A(n2252), .B(n2253), .Z(n2251) );
  CANR4CXL U2104 ( .A(n2501), .B(n1783), .C(n2699), .D(n2507), .Z(n2505) );
  CEOXL U2105 ( .A(n2513), .B(n1782), .Z(n2512) );
  CEOXL U2106 ( .A(n2227), .B(n2228), .Z(n2226) );
  CANR4CXL U2107 ( .A(n2488), .B(n1784), .C(n2690), .D(n2495), .Z(n2493) );
  CEOXL U2108 ( .A(n1783), .B(n2501), .Z(n2500) );
  CEOXL U2109 ( .A(n2201), .B(n2202), .Z(n2200) );
  CEOXL U2110 ( .A(n2214), .B(n2215), .Z(n2213) );
  CNR3XL U2111 ( .A(n2155), .B(n2657), .C(n1935), .Z(n2081) );
  CANR4CXL U2112 ( .A(n2477), .B(n1785), .C(n2691), .D(n2483), .Z(n2481) );
  CEOXL U2113 ( .A(n2488), .B(n1784), .Z(n2487) );
  CEOXL U2114 ( .A(n2175), .B(n2176), .Z(n2174) );
  CEOXL U2115 ( .A(n2188), .B(n2189), .Z(n2187) );
  CNR4XL U2116 ( .A(n2152), .B(n2153), .C(n1854), .D(n2155), .Z(n2154) );
  CANR4CXL U2117 ( .A(n2465), .B(n2656), .C(n2692), .D(n2471), .Z(n2469) );
  CEOXL U2118 ( .A(n2465), .B(n2656), .Z(n2464) );
  CEOXL U2119 ( .A(n1785), .B(n2477), .Z(n2476) );
  CANR4CXL U2120 ( .A(n2453), .B(n2452), .C(n2458), .D(n2459), .Z(n2457) );
  CEOXL U2121 ( .A(n2452), .B(n2453), .Z(n2451) );
  CNR2X1 U2122 ( .A(n2222), .B(n2677), .Z(n2233) );
  CND3X2 U2123 ( .A(n986), .B(n1890), .C(res_not_wire[26]), .Z(n2616) );
  CND3X2 U2124 ( .A(n982), .B(n1905), .C(res_not_wire[18]), .Z(n2568) );
  CND2XL U2125 ( .A(n2345), .B(n1792), .Z(n2342) );
  COND3XL U2126 ( .A(n2749), .B(n2341), .C(n2342), .D(n2343), .Z(n827) );
  CND3X2 U2127 ( .A(n987), .B(n1903), .C(res_not_wire[22]), .Z(n2592) );
  CENX1 U2128 ( .A(n102), .B(n2724), .Z(n2084) );
  COR2X1 U2129 ( .A(n2086), .B(n1937), .Z(n2724) );
  COND3XL U2130 ( .A(n2336), .B(n2748), .C(n2337), .D(n2338), .Z(n828) );
  CEOXL U2131 ( .A(res_not_wire[62]), .B(n2086), .Z(n2348) );
  COND3XL U2132 ( .A(n2749), .B(n2316), .C(n2317), .D(n2318), .Z(n831) );
  COND3XL U2133 ( .A(n2311), .B(n2748), .C(n2312), .D(n2313), .Z(n832) );
  CEOXL U2134 ( .A(res_not_wire[58]), .B(n2322), .Z(n2323) );
  CEOXL U2135 ( .A(n2309), .B(n2310), .Z(n2304) );
  COND3XL U2136 ( .A(n2748), .B(n2291), .C(n2292), .D(n2293), .Z(n835) );
  COND3XL U2137 ( .A(n2286), .B(n2747), .C(n2287), .D(n2288), .Z(n836) );
  CEOXL U2138 ( .A(n1787), .B(n2688), .Z(n2633) );
  CEOXL U2139 ( .A(res_not_wire[54]), .B(n2297), .Z(n2298) );
  CANR11XL U2140 ( .A(n1790), .B(n2641), .C(n2627), .D(n2642), .Z(n2634) );
  CEOXL U2141 ( .A(n2284), .B(n2285), .Z(n2279) );
  COND4CXL U2142 ( .A(res_not_wire[28]), .B(n1889), .C(n988), .D(n2628), .Z(
        n2622) );
  CEOXL U2143 ( .A(res_not_wire[30]), .B(n2628), .Z(n2629) );
  CEOXL U2144 ( .A(opera2[2]), .B(n1787), .Z(n2465) );
  COND3XL U2145 ( .A(n2748), .B(n2266), .C(n2267), .D(n2268), .Z(n839) );
  COND3XL U2146 ( .A(n2261), .B(n2747), .C(n2262), .D(n2263), .Z(n840) );
  CEOXL U2147 ( .A(res_not_wire[50]), .B(n2272), .Z(n2273) );
  CEOXL U2148 ( .A(n2259), .B(n2260), .Z(n2254) );
  CEOXL U2149 ( .A(n1889), .B(n1952), .Z(n2617) );
  CEOXL U2150 ( .A(opera2[4]), .B(n1787), .Z(n2477) );
  COND3XL U2151 ( .A(n2748), .B(n2241), .C(n2242), .D(n2243), .Z(n843) );
  COND4CXL U2152 ( .A(res_not_wire[26]), .B(n1890), .C(n986), .D(n2616), .Z(
        n2610) );
  CEOXL U2153 ( .A(n2234), .B(n2235), .Z(n2229) );
  CEOXL U2154 ( .A(opera2[6]), .B(n1787), .Z(n2488) );
  COND3XL U2155 ( .A(n2748), .B(n2216), .C(n2217), .D(n2218), .Z(n847) );
  COND3XL U2156 ( .A(n2236), .B(n2747), .C(n2237), .D(n2238), .Z(n844) );
  CEOXL U2157 ( .A(opera1[0]), .B(n2711), .Z(n2644) );
  CEOXL U2158 ( .A(n1891), .B(n1954), .Z(n2593) );
  CEOXL U2159 ( .A(opera2[10]), .B(n1787), .Z(n2513) );
  CEOXL U2160 ( .A(opera2[8]), .B(n1787), .Z(n2501) );
  COND3XL U2161 ( .A(n2748), .B(n2190), .C(n2191), .D(n2192), .Z(n851) );
  COND3XL U2162 ( .A(n2210), .B(n2746), .C(n2211), .D(n2212), .Z(n848) );
  CEOXL U2163 ( .A(opera1[4]), .B(n2782), .Z(n2396) );
  CEOXL U2164 ( .A(opera1[6]), .B(n2782), .Z(n2400) );
  CEOXL U2165 ( .A(opera1[3]), .B(n2782), .Z(n2394) );
  CEOXL U2166 ( .A(res_not_wire[38]), .B(n2196), .Z(n2197) );
  COND4CXL U2167 ( .A(res_not_wire[18]), .B(n1905), .C(n982), .D(n2568), .Z(
        n2562) );
  CEOXL U2168 ( .A(n1904), .B(n1956), .Z(n2569) );
  CEOXL U2169 ( .A(opera2[12]), .B(n1787), .Z(n2525) );
  CEOXL U2170 ( .A(res_not_wire[34]), .B(n1870), .Z(n2171) );
  CANR2XL U2171 ( .A(n1791), .B(result[34]), .C(result[33]), .D(n2772), .Z(
        n2161) );
  CEOXL U2172 ( .A(opera2[14]), .B(n1787), .Z(n2537) );
  CANR11XL U2173 ( .A(n2152), .B(n2153), .C(n1792), .D(n2154), .Z(n2150) );
  CANR2XL U2174 ( .A(n1791), .B(result[33]), .C(result[32]), .D(n2774), .Z(
        n2151) );
  COND4CXL U2175 ( .A(res_not_wire[8]), .B(n1922), .C(n980), .D(n2508), .Z(
        n2502) );
  COND4CXL U2176 ( .A(res_not_wire[10]), .B(n1913), .C(n979), .D(n2520), .Z(
        n2514) );
  COND4CXL U2177 ( .A(c_inres), .B(res_not_wire[0]), .C(n974), .D(n2460), .Z(
        n2454) );
  COND4CXL U2178 ( .A(res_not_wire[4]), .B(n1932), .C(n976), .D(n1927), .Z(
        n2478) );
  CEOXL U2179 ( .A(n1922), .B(n1962), .Z(n2497) );
  CEOXL U2180 ( .A(res_not_wire[2]), .B(n2460), .Z(n2461) );
  CEOXL U2181 ( .A(res_not_wire[10]), .B(n2508), .Z(n2509) );
  CEOXL U2182 ( .A(n1912), .B(n1960), .Z(n2521) );
  CEOXL U2183 ( .A(n1907), .B(n1958), .Z(n2545) );
  CEOXL U2184 ( .A(opera2[18]), .B(n1787), .Z(n2561) );
  CEOXL U2185 ( .A(opera2[16]), .B(n1787), .Z(n2549) );
  CEOXL U2186 ( .A(opera2[20]), .B(n1787), .Z(n2573) );
  CEOXL U2187 ( .A(opera2[22]), .B(n1787), .Z(n2585) );
  CEOXL U2188 ( .A(opera2[24]), .B(n1787), .Z(n2597) );
  CANR2XL U2189 ( .A(result[32]), .B(n2759), .C(n2753), .D(n1929), .Z(n2118)
         );
  CANR2XL U2190 ( .A(result[33]), .B(n2759), .C(n2753), .D(n2659), .Z(n2119)
         );
  CEOXL U2191 ( .A(opera2[26]), .B(n1787), .Z(n2609) );
  CNR2XL U2192 ( .A(n1929), .B(n2170), .Z(n2169) );
  CEOXL U2193 ( .A(opera1[26]), .B(n2777), .Z(n2440) );
  CEOXL U2194 ( .A(opera1[27]), .B(n2777), .Z(n2442) );
  CEOXL U2195 ( .A(opera2[28]), .B(n1787), .Z(n2621) );
  CEOXL U2196 ( .A(result[33]), .B(n2156), .Z(n2152) );
  CIVXL U2197 ( .A(result[32]), .Z(n1929) );
  CIVXL U2198 ( .A(res_not_wire[0]), .Z(n1968) );
  CIVXL U2199 ( .A(res_not_wire[8]), .Z(n1962) );
  CIVXL U2200 ( .A(res_not_wire[12]), .Z(n1960) );
  CIVXL U2201 ( .A(res_not_wire[16]), .Z(n1958) );
  CIVXL U2202 ( .A(res_not_wire[20]), .Z(n1956) );
  CIVXL U2203 ( .A(res_not_wire[24]), .Z(n1954) );
  CIVXL U2204 ( .A(res_not_wire[28]), .Z(n1952) );
  CND3X1 U2205 ( .A(n977), .B(n2489), .C(res_not_wire[6]), .Z(n2496) );
  CIVXL U2206 ( .A(n2489), .Z(n1927) );
  CANR4CXL U2207 ( .A(n2157), .B(n1966), .C(n2667), .D(n2163), .Z(n2162) );
  CIVX2 U2208 ( .A(n2643), .Z(n1793) );
  CNIVX1 U2209 ( .A(n1795), .Z(n2776) );
  CNIVX1 U2210 ( .A(n1795), .Z(n2772) );
  CNIVX1 U2211 ( .A(n1795), .Z(n2775) );
  CNIVX1 U2212 ( .A(n1795), .Z(n2773) );
  CNIVX1 U2213 ( .A(n1795), .Z(n2774) );
  CIVX2 U2214 ( .A(n2655), .Z(n2748) );
  CIVX2 U2215 ( .A(n2655), .Z(n2749) );
  CIVX2 U2216 ( .A(n2655), .Z(n2747) );
  CIVX2 U2217 ( .A(n2655), .Z(n2746) );
  CIVX2 U2218 ( .A(n1994), .Z(n2770) );
  CIVX2 U2219 ( .A(n2657), .Z(n2765) );
  CIVX2 U2220 ( .A(n2657), .Z(n2766) );
  CIVX2 U2221 ( .A(n2657), .Z(n2767) );
  CIVX2 U2222 ( .A(n2657), .Z(n2768) );
  CIVX2 U2223 ( .A(n2657), .Z(n2763) );
  CIVX2 U2224 ( .A(n2657), .Z(n2764) );
  CIVX2 U2225 ( .A(n2745), .Z(n2771) );
  CIVX2 U2226 ( .A(n2344), .Z(n1791) );
  CND2X1 U2227 ( .A(n1801), .B(n2082), .Z(n2643) );
  CIVX2 U2228 ( .A(n2638), .Z(n1790) );
  COND1XL U2229 ( .A(n1867), .B(n2745), .C(n1993), .Z(n2068) );
  COND1XL U2230 ( .A(n1869), .B(n1994), .C(n2743), .Z(n2058) );
  CNIVX1 U2231 ( .A(n2081), .Z(n2756) );
  CND2X1 U2232 ( .A(n1801), .B(n2743), .Z(n2745) );
  CND2X1 U2233 ( .A(n1801), .B(n2744), .Z(n1994) );
  COND1XL U2234 ( .A(n1894), .B(n1994), .C(n1993), .Z(n2038) );
  COND1XL U2235 ( .A(n1876), .B(n2745), .C(n2744), .Z(n2048) );
  CND2X1 U2236 ( .A(n2657), .B(n2071), .Z(n2744) );
  CND2X1 U2237 ( .A(n2657), .B(n2071), .Z(n2743) );
  CND2X1 U2238 ( .A(n2657), .B(n2071), .Z(n1993) );
  CNIVX1 U2239 ( .A(n2081), .Z(n2755) );
  CNIVX1 U2240 ( .A(n2081), .Z(n2754) );
  CNIVX1 U2241 ( .A(n2081), .Z(n2753) );
  CNIVX1 U2242 ( .A(n2081), .Z(n2752) );
  CNIVX1 U2243 ( .A(n2081), .Z(n2751) );
  COND2X1 U2244 ( .A(n2660), .B(n2388), .C(n2175), .D(n2176), .Z(n2182) );
  COND2X1 U2245 ( .A(n2666), .B(n2380), .C(n2227), .D(n2228), .Z(n2235) );
  COND2X1 U2246 ( .A(n2670), .B(n2375), .C(n2252), .D(n2253), .Z(n2260) );
  COND2X1 U2247 ( .A(n2675), .B(n2370), .C(n2277), .D(n2278), .Z(n2285) );
  COND2X1 U2248 ( .A(n2681), .B(n2365), .C(n2302), .D(n2303), .Z(n2310) );
  CENX1 U2249 ( .A(n2385), .B(n1980), .Z(n2195) );
  CNR3XL U2250 ( .A(n1857), .B(n2272), .C(n1943), .Z(n2283) );
  COND1XL U2251 ( .A(n1768), .B(n2398), .C(n2399), .Z(n2386) );
  CND2X1 U2252 ( .A(n2346), .B(n2347), .Z(n2355) );
  COND1XL U2253 ( .A(n2742), .B(n2352), .C(n2344), .Z(n2351) );
  CIVX2 U2254 ( .A(n2592), .Z(n1891) );
  CIVX2 U2255 ( .A(n2556), .Z(n1905) );
  CIVX2 U2256 ( .A(n2604), .Z(n1890) );
  CIVX2 U2257 ( .A(n2580), .Z(n1903) );
  CENX1 U2258 ( .A(n2381), .B(n1978), .Z(n2220) );
  CENX1 U2259 ( .A(n2376), .B(n1976), .Z(n2245) );
  CENX1 U2260 ( .A(n2371), .B(n1974), .Z(n2270) );
  CENX1 U2261 ( .A(n2366), .B(n1972), .Z(n2295) );
  COND1XL U2262 ( .A(n1760), .B(n2412), .C(n2413), .Z(n2379) );
  COND1XL U2263 ( .A(n1754), .B(n2420), .C(n2421), .Z(n2374) );
  COND1XL U2264 ( .A(n1748), .B(n2428), .C(n2429), .Z(n2369) );
  COND1XL U2265 ( .A(n1764), .B(n2406), .C(n2407), .Z(n2382) );
  COND1XL U2266 ( .A(n1758), .B(n2414), .C(n2415), .Z(n2377) );
  COND1XL U2267 ( .A(n1752), .B(n2422), .C(n2423), .Z(n2372) );
  COND1XL U2268 ( .A(n1766), .B(n2402), .C(n2403), .Z(n2384) );
  COND1XL U2269 ( .A(n1762), .B(n2410), .C(n2411), .Z(n2380) );
  COND1XL U2270 ( .A(n1756), .B(n2418), .C(n2419), .Z(n2375) );
  COND1XL U2271 ( .A(n1750), .B(n2426), .C(n2427), .Z(n2370) );
  CND2X1 U2272 ( .A(n1762), .B(n2410), .Z(n2411) );
  CND2X1 U2273 ( .A(n1760), .B(n2412), .Z(n2413) );
  CND2X1 U2274 ( .A(n1758), .B(n2414), .Z(n2415) );
  CND2X1 U2275 ( .A(n1756), .B(n2418), .Z(n2419) );
  CND2X1 U2276 ( .A(n1754), .B(n2420), .Z(n2421) );
  CND2X1 U2277 ( .A(n1752), .B(n2422), .Z(n2423) );
  CND2X1 U2278 ( .A(n1750), .B(n2426), .Z(n2427) );
  CND2X1 U2279 ( .A(n1748), .B(n2428), .Z(n2429) );
  CND2X1 U2280 ( .A(n1746), .B(n2430), .Z(n2431) );
  CND2X1 U2281 ( .A(n1757), .B(n2416), .Z(n2417) );
  CND2X1 U2282 ( .A(n1751), .B(n2424), .Z(n2425) );
  CND2X1 U2283 ( .A(n1745), .B(n2432), .Z(n2433) );
  CENX1 U2284 ( .A(n2361), .B(n1970), .Z(n2320) );
  COND1XL U2285 ( .A(n1742), .B(n2436), .C(n2437), .Z(n2364) );
  COND1XL U2286 ( .A(n1736), .B(n2444), .C(n2445), .Z(n2359) );
  COND1XL U2287 ( .A(n1746), .B(n2430), .C(n2431), .Z(n2367) );
  COND1XL U2288 ( .A(n1740), .B(n2438), .C(n2439), .Z(n2362) );
  COND1XL U2289 ( .A(n1734), .B(n2446), .C(n2354), .Z(n2357) );
  COND1XL U2290 ( .A(n1744), .B(n2434), .C(n2435), .Z(n2365) );
  COND1XL U2291 ( .A(n1738), .B(n2442), .C(n2443), .Z(n2360) );
  CENX1 U2292 ( .A(n2447), .B(n2353), .Z(n2346) );
  CEOX1 U2293 ( .A(n2354), .B(n1983), .Z(n2447) );
  CND2X1 U2294 ( .A(n1734), .B(n2446), .Z(n2354) );
  CND2X1 U2295 ( .A(n1744), .B(n2434), .Z(n2435) );
  CND2X1 U2296 ( .A(n1742), .B(n2436), .Z(n2437) );
  CND2X1 U2297 ( .A(n1740), .B(n2438), .Z(n2439) );
  CND2X1 U2298 ( .A(n1738), .B(n2442), .Z(n2443) );
  CND2X1 U2299 ( .A(n1736), .B(n2444), .Z(n2445) );
  CND2X1 U2300 ( .A(n1739), .B(n2440), .Z(n2441) );
  COND3X1 U2301 ( .A(n1995), .B(n2071), .C(n2076), .D(n2645), .Z(n2082) );
  CND2X1 U2302 ( .A(n1793), .B(n1854), .Z(n2344) );
  CNR3XL U2303 ( .A(n1986), .B(n1985), .C(n1930), .Z(n1999) );
  CIVX2 U2304 ( .A(n2742), .Z(n1792) );
  CND2X1 U2305 ( .A(n1990), .B(n2082), .Z(n2638) );
  COND2X1 U2306 ( .A(n2051), .B(n1878), .C(n1994), .D(n2052), .Z(n931) );
  CND2X1 U2307 ( .A(n1875), .B(n1878), .Z(n2052) );
  COND2X1 U2308 ( .A(n2061), .B(n1872), .C(n2745), .D(n2062), .Z(n927) );
  CND2X1 U2309 ( .A(n1868), .B(n1872), .Z(n2062) );
  CNIVX1 U2310 ( .A(n2080), .Z(n2762) );
  COND2X1 U2311 ( .A(n1880), .B(n2744), .C(n1866), .D(n2745), .Z(n955) );
  CANR1XL U2312 ( .A(n1797), .B(n1990), .C(n2078), .Z(n2645) );
  CND3XL U2313 ( .A(n2073), .B(n2076), .C(n2077), .Z(n1989) );
  CANR3X1 U2314 ( .A(n1936), .B(n1803), .C(n2078), .D(n1800), .Z(n2077) );
  CNIVX1 U2315 ( .A(n2080), .Z(n2758) );
  CNIVX1 U2316 ( .A(n2080), .Z(n2757) );
  CND2X1 U2317 ( .A(n1801), .B(n2646), .Z(n2071) );
  COND2X1 U2318 ( .A(n2021), .B(n1920), .C(n1994), .D(n2022), .Z(n943) );
  CND2X1 U2319 ( .A(n2023), .B(n1920), .Z(n2022) );
  COND2X1 U2320 ( .A(n2011), .B(n1917), .C(n1994), .D(n2012), .Z(n947) );
  CND2X1 U2321 ( .A(n2013), .B(n1917), .Z(n2012) );
  COND2X1 U2322 ( .A(n2016), .B(n1916), .C(n2745), .D(n2017), .Z(n945) );
  CND2X1 U2323 ( .A(n2018), .B(n1916), .Z(n2017) );
  COND2X1 U2324 ( .A(n2026), .B(n1901), .C(n2745), .D(n2027), .Z(n941) );
  CND2X1 U2325 ( .A(n2028), .B(n1901), .Z(n2027) );
  COND2X1 U2326 ( .A(n2031), .B(n1899), .C(n1994), .D(n2032), .Z(n939) );
  CND2X1 U2327 ( .A(n1898), .B(n1899), .Z(n2032) );
  COND2X1 U2328 ( .A(n2041), .B(n1893), .C(n2745), .D(n2042), .Z(n935) );
  CND2X1 U2329 ( .A(n1884), .B(n1893), .Z(n2042) );
  COND3X1 U2330 ( .A(n2000), .B(n1926), .C(n2001), .D(n1998), .Z(n953) );
  CND3XL U2331 ( .A(n2002), .B(n1926), .C(n2770), .Z(n2001) );
  COND3X1 U2332 ( .A(n1996), .B(n1925), .C(n1997), .D(n1998), .Z(n954) );
  CND3XL U2333 ( .A(n1999), .B(n1925), .C(n2770), .Z(n1997) );
  CNIVX1 U2334 ( .A(n2080), .Z(n2761) );
  CNIVX1 U2335 ( .A(n2080), .Z(n2760) );
  CNIVX1 U2336 ( .A(n2080), .Z(n2759) );
  COND3X1 U2337 ( .A(n1989), .B(n1819), .C(n2074), .D(n2075), .Z(n921) );
  CND2X1 U2338 ( .A(n1988), .B(n1989), .Z(n2074) );
  CND3XL U2339 ( .A(n1895), .B(n1893), .C(n1920), .Z(n2648) );
  CNR2IX1 U2340 ( .B(n2071), .A(n1990), .Z(n2073) );
  COND1XL U2341 ( .A(n1989), .B(n2708), .C(n2073), .Z(n922) );
  CANR2X1 U2342 ( .A(n2391), .B(n2659), .C(n1770), .D(n2153), .Z(n2390) );
  CANR2X1 U2343 ( .A(result[36]), .B(n2387), .C(n2182), .D(n2183), .Z(n2188)
         );
  CANR2X1 U2344 ( .A(result[42]), .B(n2381), .C(n2221), .D(n2220), .Z(n2227)
         );
  CEOX1 U2345 ( .A(n2387), .B(result[36]), .Z(n2183) );
  CEOX1 U2346 ( .A(result[37]), .B(n2386), .Z(n2189) );
  CEOX1 U2347 ( .A(result[35]), .B(n2388), .Z(n2176) );
  CNR3XL U2348 ( .A(n2297), .B(n110), .C(n1941), .Z(n2308) );
  CEOX1 U2349 ( .A(n2383), .B(result[40]), .Z(n2209) );
  CANR2X1 U2350 ( .A(result[40]), .B(n2383), .C(n2208), .D(n2209), .Z(n2214)
         );
  CANR2X1 U2351 ( .A(result[38]), .B(n2385), .C(n2194), .D(n2195), .Z(n2201)
         );
  CANR2X1 U2352 ( .A(result[46]), .B(n2376), .C(n2246), .D(n2245), .Z(n2252)
         );
  CANR2X1 U2353 ( .A(result[50]), .B(n2371), .C(n2271), .D(n2270), .Z(n2277)
         );
  CANR2X1 U2354 ( .A(result[54]), .B(n2366), .C(n2296), .D(n2295), .Z(n2302)
         );
  CANR2X1 U2355 ( .A(result[58]), .B(n2361), .C(n2321), .D(n2320), .Z(n2327)
         );
  CNR3XL U2356 ( .A(n2322), .B(n106), .C(n1939), .Z(n2333) );
  COND1XL U2357 ( .A(c_inop1), .B(n2644), .C(n2393), .Z(n2170) );
  COND2X1 U2358 ( .A(n2082), .B(n1851), .C(n2750), .D(n2084), .Z(n919) );
  CND2X1 U2359 ( .A(n1772), .B(result[32]), .Z(n2153) );
  COND3X1 U2360 ( .A(n2742), .B(n2329), .C(n2330), .D(n2331), .Z(n829) );
  CANR2X1 U2361 ( .A(n1791), .B(result[60]), .C(result[59]), .D(n2774), .Z(
        n2331) );
  CND2X1 U2362 ( .A(n2332), .B(n2655), .Z(n2330) );
  CANR2X1 U2363 ( .A(n1791), .B(result[62]), .C(result[61]), .D(n2774), .Z(
        n2343) );
  COND3X1 U2364 ( .A(n2348), .B(n2748), .C(n2349), .D(n2350), .Z(n826) );
  CND3XL U2365 ( .A(n2352), .B(n1851), .C(n1792), .Z(n2349) );
  CANR2X1 U2366 ( .A(result[63]), .B(n2351), .C(result[62]), .D(n2774), .Z(
        n2350) );
  CANR2X1 U2367 ( .A(n1791), .B(result[61]), .C(result[60]), .D(n2774), .Z(
        n2338) );
  CND2X1 U2368 ( .A(n2339), .B(n1792), .Z(n2337) );
  CEOX1 U2369 ( .A(n2379), .B(result[44]), .Z(n2234) );
  CEOX1 U2370 ( .A(n2374), .B(result[48]), .Z(n2259) );
  CEOX1 U2371 ( .A(n2369), .B(result[52]), .Z(n2284) );
  CEOX1 U2372 ( .A(result[41]), .B(n2382), .Z(n2215) );
  CEOX1 U2373 ( .A(result[45]), .B(n2377), .Z(n2240) );
  CEOX1 U2374 ( .A(result[49]), .B(n2372), .Z(n2265) );
  CEOX1 U2375 ( .A(result[39]), .B(n2384), .Z(n2202) );
  CEOX1 U2376 ( .A(result[43]), .B(n2380), .Z(n2228) );
  CEOX1 U2377 ( .A(result[47]), .B(n2375), .Z(n2253) );
  CEOX1 U2378 ( .A(result[51]), .B(n2370), .Z(n2278) );
  COND4CX1 U2379 ( .A(res_not_wire[30]), .B(n1883), .C(n989), .D(n2157), .Z(
        n2637) );
  CEOX1 U2380 ( .A(n2704), .B(opera2[31]), .Z(n2640) );
  CEOX1 U2381 ( .A(opera1[5]), .B(n2781), .Z(n2398) );
  COND3X1 U2382 ( .A(n2742), .B(n2279), .C(n2280), .D(n2281), .Z(n837) );
  CANR2X1 U2383 ( .A(n1791), .B(result[52]), .C(result[51]), .D(n2773), .Z(
        n2281) );
  CND2X1 U2384 ( .A(n2282), .B(n2655), .Z(n2280) );
  CANR2X1 U2385 ( .A(n1791), .B(result[54]), .C(result[53]), .D(n2773), .Z(
        n2293) );
  CND2X1 U2386 ( .A(n2294), .B(n1792), .Z(n2292) );
  COND3X1 U2387 ( .A(n2742), .B(n2304), .C(n2305), .D(n2306), .Z(n833) );
  CANR2X1 U2388 ( .A(n1791), .B(result[56]), .C(result[55]), .D(n2773), .Z(
        n2306) );
  CND2X1 U2389 ( .A(n2307), .B(n2655), .Z(n2305) );
  CANR2X1 U2390 ( .A(n1791), .B(result[58]), .C(result[57]), .D(n2773), .Z(
        n2318) );
  CND2X1 U2391 ( .A(n2319), .B(n1792), .Z(n2317) );
  CANR2X1 U2392 ( .A(n1791), .B(result[53]), .C(result[52]), .D(n2773), .Z(
        n2288) );
  CND2X1 U2393 ( .A(n2289), .B(n1792), .Z(n2287) );
  COND3X1 U2394 ( .A(n2298), .B(n2748), .C(n2299), .D(n2300), .Z(n834) );
  CANR2X1 U2395 ( .A(n1791), .B(result[55]), .C(result[54]), .D(n2773), .Z(
        n2300) );
  CND2X1 U2396 ( .A(n2301), .B(n1792), .Z(n2299) );
  CANR2X1 U2397 ( .A(n1791), .B(result[57]), .C(result[56]), .D(n2773), .Z(
        n2313) );
  CND2X1 U2398 ( .A(n2314), .B(n1792), .Z(n2312) );
  COND3X1 U2399 ( .A(n2323), .B(n2748), .C(n2324), .D(n2325), .Z(n830) );
  CANR2X1 U2400 ( .A(n1791), .B(result[59]), .C(result[58]), .D(n2774), .Z(
        n2325) );
  CND2X1 U2401 ( .A(n2326), .B(n1792), .Z(n2324) );
  COND3X1 U2402 ( .A(n2629), .B(n2746), .C(n2630), .D(n2631), .Z(n795) );
  CANR2X1 U2403 ( .A(n1793), .B(result[31]), .C(result[30]), .D(n2772), .Z(
        n2631) );
  CND2X1 U2404 ( .A(n1790), .B(n2632), .Z(n2630) );
  CEOX1 U2405 ( .A(n2364), .B(result[56]), .Z(n2309) );
  CEOX1 U2406 ( .A(result[53]), .B(n2367), .Z(n2290) );
  CEOX1 U2407 ( .A(result[57]), .B(n2362), .Z(n2315) );
  CEOX1 U2408 ( .A(result[61]), .B(n2357), .Z(n2340) );
  CEOX1 U2409 ( .A(result[55]), .B(n2365), .Z(n2303) );
  CEOX1 U2410 ( .A(result[59]), .B(n2360), .Z(n2328) );
  CENX1 U2411 ( .A(opera1[2]), .B(n2783), .Z(n2167) );
  CEOX1 U2412 ( .A(opera1[7]), .B(n2781), .Z(n2402) );
  CEOX1 U2413 ( .A(opera1[9]), .B(n2781), .Z(n2406) );
  CEOX1 U2414 ( .A(n2359), .B(result[60]), .Z(n2334) );
  CEOX1 U2415 ( .A(opera1[8]), .B(n2781), .Z(n2404) );
  CEOX1 U2416 ( .A(opera1[10]), .B(n2781), .Z(n2408) );
  COND3X1 U2417 ( .A(n2742), .B(n2229), .C(n2230), .D(n2231), .Z(n845) );
  CANR2X1 U2418 ( .A(n1791), .B(result[44]), .C(result[43]), .D(n2772), .Z(
        n2231) );
  CND2X1 U2419 ( .A(n2232), .B(n2655), .Z(n2230) );
  CANR2X1 U2420 ( .A(n1791), .B(result[46]), .C(result[45]), .D(n2773), .Z(
        n2243) );
  CND2X1 U2421 ( .A(n2244), .B(n1792), .Z(n2242) );
  COND3X1 U2422 ( .A(n2742), .B(n2254), .C(n2255), .D(n2256), .Z(n841) );
  CANR2X1 U2423 ( .A(n1791), .B(result[48]), .C(result[47]), .D(n2773), .Z(
        n2256) );
  CND2X1 U2424 ( .A(n2257), .B(n2655), .Z(n2255) );
  CANR2X1 U2425 ( .A(n1791), .B(result[50]), .C(result[49]), .D(n2774), .Z(
        n2268) );
  CND2X1 U2426 ( .A(n2269), .B(n1792), .Z(n2267) );
  CND2X1 U2427 ( .A(n2239), .B(n1792), .Z(n2237) );
  CANR2X1 U2428 ( .A(n1791), .B(result[45]), .C(result[44]), .D(n2772), .Z(
        n2238) );
  COND3X1 U2429 ( .A(n2248), .B(n2747), .C(n2249), .D(n2250), .Z(n842) );
  CND2X1 U2430 ( .A(n2251), .B(n1792), .Z(n2249) );
  CANR2X1 U2431 ( .A(n1791), .B(result[47]), .C(result[46]), .D(n2773), .Z(
        n2250) );
  CEOX1 U2432 ( .A(res_not_wire[46]), .B(n2247), .Z(n2248) );
  CANR2X1 U2433 ( .A(n1791), .B(result[49]), .C(result[48]), .D(n2773), .Z(
        n2263) );
  CND2X1 U2434 ( .A(n2264), .B(n1792), .Z(n2262) );
  COND3X1 U2435 ( .A(n2273), .B(n2747), .C(n2274), .D(n2275), .Z(n838) );
  CANR2X1 U2436 ( .A(n1791), .B(result[51]), .C(result[50]), .D(n2773), .Z(
        n2275) );
  CND2X1 U2437 ( .A(n2276), .B(n1792), .Z(n2274) );
  COND3X1 U2438 ( .A(n2750), .B(n2610), .C(n2611), .D(n2612), .Z(n798) );
  CANR2X1 U2439 ( .A(n1793), .B(result[28]), .C(result[27]), .D(n2776), .Z(
        n2612) );
  CND2X1 U2440 ( .A(n2613), .B(n1790), .Z(n2611) );
  COND3X1 U2441 ( .A(n2750), .B(n2622), .C(n2623), .D(n2624), .Z(n796) );
  CANR2X1 U2442 ( .A(n1793), .B(result[30]), .C(result[29]), .D(n2776), .Z(
        n2624) );
  CND2X1 U2443 ( .A(n2625), .B(n1790), .Z(n2623) );
  COND3X1 U2444 ( .A(n2605), .B(n2746), .C(n2606), .D(n2607), .Z(n799) );
  CANR2X1 U2445 ( .A(n1793), .B(result[27]), .C(result[26]), .D(n2776), .Z(
        n2607) );
  CND2X1 U2446 ( .A(n1790), .B(n2608), .Z(n2606) );
  CANR2X1 U2447 ( .A(n1793), .B(result[29]), .C(result[28]), .D(n2776), .Z(
        n2619) );
  CND2X1 U2448 ( .A(n1790), .B(n2620), .Z(n2618) );
  CEOX1 U2449 ( .A(opera1[11]), .B(n2780), .Z(n2410) );
  CEOX1 U2450 ( .A(opera1[12]), .B(n2780), .Z(n2412) );
  CEOX1 U2451 ( .A(opera1[13]), .B(n2780), .Z(n2414) );
  CEOX1 U2452 ( .A(opera1[14]), .B(n2780), .Z(n2416) );
  CND2X1 U2453 ( .A(n2193), .B(n1792), .Z(n2191) );
  CANR2X1 U2454 ( .A(n1791), .B(result[38]), .C(result[37]), .D(n2772), .Z(
        n2192) );
  CND2X1 U2455 ( .A(n2219), .B(n1792), .Z(n2217) );
  CANR2X1 U2456 ( .A(n1791), .B(result[42]), .C(result[41]), .D(n2772), .Z(
        n2218) );
  COND3X1 U2457 ( .A(n2184), .B(n2746), .C(n2185), .D(n2186), .Z(n852) );
  CND2X1 U2458 ( .A(n2187), .B(n1792), .Z(n2185) );
  CANR2X1 U2459 ( .A(n1791), .B(result[37]), .C(result[36]), .D(n2773), .Z(
        n2186) );
  COND3X1 U2460 ( .A(n2197), .B(n2746), .C(n2198), .D(n2199), .Z(n850) );
  CND2X1 U2461 ( .A(n2200), .B(n1792), .Z(n2198) );
  CANR2X1 U2462 ( .A(n1791), .B(result[39]), .C(result[38]), .D(n2772), .Z(
        n2199) );
  CND2X1 U2463 ( .A(n2213), .B(n1792), .Z(n2211) );
  CANR2X1 U2464 ( .A(n1791), .B(result[41]), .C(result[40]), .D(n2772), .Z(
        n2212) );
  COND3X1 U2465 ( .A(n2223), .B(n2746), .C(n2224), .D(n2225), .Z(n846) );
  CND2X1 U2466 ( .A(n2226), .B(n1792), .Z(n2224) );
  CANR2X1 U2467 ( .A(n1791), .B(result[43]), .C(result[42]), .D(n2772), .Z(
        n2225) );
  CEOX1 U2468 ( .A(res_not_wire[42]), .B(n2222), .Z(n2223) );
  COND3X1 U2469 ( .A(n2750), .B(n2586), .C(n2587), .D(n2588), .Z(n802) );
  CANR2X1 U2470 ( .A(n1793), .B(result[24]), .C(result[23]), .D(n2776), .Z(
        n2588) );
  CND2X1 U2471 ( .A(n2589), .B(n1790), .Z(n2587) );
  COND3X1 U2472 ( .A(n2750), .B(n2598), .C(n2599), .D(n2600), .Z(n800) );
  CANR2X1 U2473 ( .A(n1793), .B(result[26]), .C(result[25]), .D(n2776), .Z(
        n2600) );
  CND2X1 U2474 ( .A(n2601), .B(n1790), .Z(n2599) );
  CANR2X1 U2475 ( .A(n1793), .B(result[25]), .C(result[24]), .D(n2776), .Z(
        n2595) );
  CND2X1 U2476 ( .A(n1790), .B(n2596), .Z(n2594) );
  COND3X1 U2477 ( .A(n2742), .B(n2177), .C(n2178), .D(n2179), .Z(n853) );
  CENX1 U2478 ( .A(n2182), .B(n2183), .Z(n2177) );
  CANR2X1 U2479 ( .A(n1791), .B(result[36]), .C(result[35]), .D(n2772), .Z(
        n2179) );
  CND2X1 U2480 ( .A(n2180), .B(n2655), .Z(n2178) );
  COND3X1 U2481 ( .A(n2742), .B(n2203), .C(n2204), .D(n2205), .Z(n849) );
  CANR2X1 U2482 ( .A(n1791), .B(result[40]), .C(result[39]), .D(n2772), .Z(
        n2205) );
  CND2X1 U2483 ( .A(n2206), .B(n2655), .Z(n2204) );
  CANR11X1 U2484 ( .A(i[30]), .B(n1867), .C(i[29]), .D(n1880), .Z(n1995) );
  COND3X1 U2485 ( .A(n2149), .B(n2746), .C(n2150), .D(n2151), .Z(n856) );
  CEOX1 U2486 ( .A(n2157), .B(res_not_wire[32]), .Z(n2149) );
  COND3X1 U2487 ( .A(n2448), .B(n2748), .C(n2449), .D(n2450), .Z(n825) );
  CEOX1 U2488 ( .A(n1968), .B(c_inres), .Z(n2448) );
  CND2X1 U2489 ( .A(n1790), .B(n2451), .Z(n2449) );
  CANR2X1 U2490 ( .A(n1793), .B(result[1]), .C(n2772), .D(result[0]), .Z(n2450) );
  COND3X1 U2491 ( .A(n2749), .B(n2502), .C(n2503), .D(n2504), .Z(n816) );
  CND2X1 U2492 ( .A(n2505), .B(n1790), .Z(n2503) );
  CANR2X1 U2493 ( .A(n1793), .B(result[10]), .C(result[9]), .D(n2775), .Z(
        n2504) );
  COND3X1 U2494 ( .A(n2749), .B(n2514), .C(n2515), .D(n2516), .Z(n814) );
  CND2X1 U2495 ( .A(n2517), .B(n1790), .Z(n2515) );
  CANR2X1 U2496 ( .A(n1793), .B(result[12]), .C(result[11]), .D(n2775), .Z(
        n2516) );
  COND3X1 U2497 ( .A(n2749), .B(n2526), .C(n2527), .D(n2528), .Z(n812) );
  CND2X1 U2498 ( .A(n2529), .B(n1790), .Z(n2527) );
  CANR2X1 U2499 ( .A(n1793), .B(result[14]), .C(result[13]), .D(n2775), .Z(
        n2528) );
  COND3X1 U2500 ( .A(n2749), .B(n2538), .C(n2539), .D(n2540), .Z(n810) );
  CND2X1 U2501 ( .A(n2541), .B(n1790), .Z(n2539) );
  CANR2X1 U2502 ( .A(n1793), .B(result[16]), .C(result[15]), .D(n2775), .Z(
        n2540) );
  COND3X1 U2503 ( .A(n2749), .B(n2550), .C(n2551), .D(n2552), .Z(n808) );
  CND2X1 U2504 ( .A(n2553), .B(n1790), .Z(n2551) );
  CANR2X1 U2505 ( .A(n1793), .B(result[18]), .C(result[17]), .D(n2775), .Z(
        n2552) );
  COND3X1 U2506 ( .A(n2749), .B(n2562), .C(n2563), .D(n2564), .Z(n806) );
  CND2X1 U2507 ( .A(n2565), .B(n1790), .Z(n2563) );
  CANR2X1 U2508 ( .A(n1793), .B(result[20]), .C(result[19]), .D(n2775), .Z(
        n2564) );
  COND3X1 U2509 ( .A(n2749), .B(n2454), .C(n2455), .D(n2456), .Z(n824) );
  CND2X1 U2510 ( .A(n2457), .B(n1790), .Z(n2455) );
  CANR2X1 U2511 ( .A(n1793), .B(result[2]), .C(result[1]), .D(n2774), .Z(n2456) );
  COND3X1 U2512 ( .A(n2749), .B(n2466), .C(n2467), .D(n2468), .Z(n822) );
  CND2X1 U2513 ( .A(n2469), .B(n1790), .Z(n2467) );
  CANR2X1 U2514 ( .A(n1793), .B(result[4]), .C(result[3]), .D(n2774), .Z(n2468) );
  COND3X1 U2515 ( .A(n2749), .B(n2478), .C(n2479), .D(n2480), .Z(n820) );
  CND2X1 U2516 ( .A(n2481), .B(n1790), .Z(n2479) );
  CANR2X1 U2517 ( .A(n1793), .B(result[6]), .C(result[5]), .D(n2774), .Z(n2480) );
  COND3X1 U2518 ( .A(n2749), .B(n2490), .C(n2491), .D(n2492), .Z(n818) );
  CND2X1 U2519 ( .A(n2493), .B(n1790), .Z(n2491) );
  CANR2X1 U2520 ( .A(n1793), .B(result[8]), .C(result[7]), .D(n2775), .Z(n2492) );
  CND2X1 U2521 ( .A(n1790), .B(n2500), .Z(n2498) );
  CANR2X1 U2522 ( .A(n1793), .B(result[9]), .C(result[8]), .D(n2775), .Z(n2499) );
  COND3X1 U2523 ( .A(n2461), .B(n2748), .C(n2462), .D(n2463), .Z(n823) );
  CND2X1 U2524 ( .A(n1790), .B(n2464), .Z(n2462) );
  CANR2X1 U2525 ( .A(n1793), .B(result[3]), .C(result[2]), .D(n2774), .Z(n2463) );
  CND2X1 U2526 ( .A(n1790), .B(n2476), .Z(n2474) );
  CANR2X1 U2527 ( .A(n1793), .B(result[5]), .C(result[4]), .D(n2774), .Z(n2475) );
  COND3X1 U2528 ( .A(n2484), .B(n2747), .C(n2485), .D(n2486), .Z(n819) );
  CEOX1 U2529 ( .A(res_not_wire[6]), .B(n1927), .Z(n2484) );
  CND2X1 U2530 ( .A(n1790), .B(n2487), .Z(n2485) );
  CANR2X1 U2531 ( .A(n1793), .B(result[7]), .C(result[6]), .D(n2774), .Z(n2486) );
  COND3X1 U2532 ( .A(n2509), .B(n2747), .C(n2510), .D(n2511), .Z(n815) );
  CND2X1 U2533 ( .A(n1790), .B(n2512), .Z(n2510) );
  CANR2X1 U2534 ( .A(n1793), .B(result[11]), .C(result[10]), .D(n2775), .Z(
        n2511) );
  COND3X1 U2535 ( .A(n2521), .B(n2747), .C(n2522), .D(n2523), .Z(n813) );
  CND2X1 U2536 ( .A(n1790), .B(n2524), .Z(n2522) );
  CANR2X1 U2537 ( .A(n1793), .B(result[13]), .C(result[12]), .D(n2775), .Z(
        n2523) );
  COND3X1 U2538 ( .A(n2533), .B(n2747), .C(n2534), .D(n2535), .Z(n811) );
  CND2X1 U2539 ( .A(n1790), .B(n2536), .Z(n2534) );
  CANR2X1 U2540 ( .A(n1793), .B(result[15]), .C(result[14]), .D(n2775), .Z(
        n2535) );
  COND3X1 U2541 ( .A(n2545), .B(n2747), .C(n2546), .D(n2547), .Z(n809) );
  CND2X1 U2542 ( .A(n1790), .B(n2548), .Z(n2546) );
  CANR2X1 U2543 ( .A(n1793), .B(result[17]), .C(result[16]), .D(n2775), .Z(
        n2547) );
  COND3X1 U2544 ( .A(n2557), .B(n2747), .C(n2558), .D(n2559), .Z(n807) );
  CND2X1 U2545 ( .A(n1790), .B(n2560), .Z(n2558) );
  CANR2X1 U2546 ( .A(n1793), .B(result[19]), .C(result[18]), .D(n2775), .Z(
        n2559) );
  CEOX1 U2547 ( .A(opera1[15]), .B(n2779), .Z(n2418) );
  CEOX1 U2548 ( .A(opera1[16]), .B(n2779), .Z(n2420) );
  CEOX1 U2549 ( .A(opera1[17]), .B(n2779), .Z(n2422) );
  CEOX1 U2550 ( .A(opera1[18]), .B(n2779), .Z(n2424) );
  CND3XL U2551 ( .A(i[23]), .B(n1875), .C(i[24]), .Z(n2056) );
  CND3XL U2552 ( .A(i[19]), .B(n1884), .C(i[20]), .Z(n2046) );
  CND3XL U2553 ( .A(i[27]), .B(n1868), .C(i[28]), .Z(n2066) );
  COND3X1 U2554 ( .A(n2158), .B(n2742), .C(n2160), .D(n2161), .Z(n855) );
  CEOX1 U2555 ( .A(n2164), .B(n2165), .Z(n2158) );
  CND2X1 U2556 ( .A(n2162), .B(n2655), .Z(n2160) );
  COND3X1 U2557 ( .A(n2171), .B(n2746), .C(n2172), .D(n2173), .Z(n854) );
  CND2X1 U2558 ( .A(n2174), .B(n1792), .Z(n2172) );
  CANR2X1 U2559 ( .A(n1791), .B(result[35]), .C(result[34]), .D(n2772), .Z(
        n2173) );
  CND3XL U2560 ( .A(i[15]), .B(n1898), .C(i[16]), .Z(n2036) );
  CND3XL U2561 ( .A(i[13]), .B(n2028), .C(i[14]), .Z(n2035) );
  CND3XL U2562 ( .A(i[17]), .B(n1894), .C(i[18]), .Z(n2045) );
  CND3XL U2563 ( .A(i[25]), .B(n1869), .C(i[26]), .Z(n2065) );
  CND3XL U2564 ( .A(i[21]), .B(n1876), .C(i[22]), .Z(n2055) );
  COND3X1 U2565 ( .A(n2749), .B(n2574), .C(n2575), .D(n2576), .Z(n804) );
  CANR2X1 U2566 ( .A(n1793), .B(result[22]), .C(result[21]), .D(n2776), .Z(
        n2576) );
  CND2X1 U2567 ( .A(n2577), .B(n1790), .Z(n2575) );
  CANR2X1 U2568 ( .A(n1793), .B(result[21]), .C(result[20]), .D(n2776), .Z(
        n2571) );
  CND2X1 U2569 ( .A(n1790), .B(n2572), .Z(n2570) );
  COND3X1 U2570 ( .A(n2581), .B(n2746), .C(n2582), .D(n2583), .Z(n803) );
  CANR2X1 U2571 ( .A(n1793), .B(result[23]), .C(result[22]), .D(n2776), .Z(
        n2583) );
  CND2X1 U2572 ( .A(n1790), .B(n2584), .Z(n2582) );
  CNIVX1 U2573 ( .A(n2159), .Z(n2742) );
  CND2X1 U2574 ( .A(n1793), .B(result[0]), .Z(n2159) );
  CEOX1 U2575 ( .A(opera1[19]), .B(n2779), .Z(n2426) );
  CEOX1 U2576 ( .A(opera1[20]), .B(n2778), .Z(n2428) );
  CEOX1 U2577 ( .A(opera1[21]), .B(n2778), .Z(n2430) );
  CNR3XL U2578 ( .A(n2657), .B(n1007), .C(n2155), .Z(n2080) );
  CND3XL U2579 ( .A(n1925), .B(n1923), .C(n1930), .Z(n2651) );
  CEOX1 U2580 ( .A(opera1[23]), .B(n2778), .Z(n2434) );
  CEOX1 U2581 ( .A(opera1[24]), .B(n2780), .Z(n2436) );
  CEOX1 U2582 ( .A(opera1[25]), .B(n2778), .Z(n2438) );
  COND11X1 U2583 ( .A(n2745), .B(i[29]), .C(n2066), .D(n2067), .Z(n925) );
  CND2X1 U2584 ( .A(i[29]), .B(n2068), .Z(n2067) );
  COND11X1 U2585 ( .A(n1994), .B(i[25]), .C(n2056), .D(n2057), .Z(n929) );
  CND2X1 U2586 ( .A(i[25]), .B(n2058), .Z(n2057) );
  CEOX1 U2587 ( .A(opera1[22]), .B(n2778), .Z(n2432) );
  CND4X1 U2588 ( .A(n1887), .B(n1924), .C(n1917), .D(n1915), .Z(n2654) );
  CND4X1 U2589 ( .A(n1900), .B(n1899), .C(n1885), .D(n1878), .Z(n2653) );
  COND1XL U2590 ( .A(n2763), .B(n1933), .C(n2087), .Z(n918) );
  CANR2X1 U2591 ( .A(result[1]), .B(n2762), .C(n2756), .D(n1840), .Z(n2087) );
  COND1XL U2592 ( .A(n2763), .B(n1931), .C(n2089), .Z(n916) );
  CANR2X1 U2593 ( .A(result[3]), .B(n2762), .C(n2756), .D(n1839), .Z(n2089) );
  COND1XL U2594 ( .A(n2763), .B(n1968), .C(n2079), .Z(n920) );
  CANR2X1 U2595 ( .A(result[0]), .B(n2762), .C(n2756), .D(n1854), .Z(n2079) );
  COND1XL U2596 ( .A(n2763), .B(n1965), .C(n2088), .Z(n917) );
  CANR2X1 U2597 ( .A(result[2]), .B(n2762), .C(n2756), .D(n1834), .Z(n2088) );
  COND4CX1 U2598 ( .A(n2061), .B(n2063), .C(n1873), .D(n2064), .Z(n926) );
  CND2X1 U2599 ( .A(n2770), .B(n1872), .Z(n2063) );
  COND4CX1 U2600 ( .A(n2051), .B(n2053), .C(n1865), .D(n2054), .Z(n930) );
  CND2X1 U2601 ( .A(n2770), .B(n1878), .Z(n2053) );
  CND2X1 U2602 ( .A(n1880), .B(n2652), .Z(n2646) );
  CND2X1 U2603 ( .A(n2059), .B(n2060), .Z(n928) );
  COND4CX1 U2604 ( .A(n2770), .B(n1877), .C(n2058), .D(i[26]), .Z(n2059) );
  CND2X1 U2605 ( .A(n2069), .B(n2070), .Z(n924) );
  COND4CX1 U2606 ( .A(n2770), .B(n1887), .C(n2068), .D(i[30]), .Z(n2069) );
  CNR3XL U2607 ( .A(n1936), .B(n56), .C(n1803), .Z(n1990) );
  CND3XL U2608 ( .A(n1368), .B(n1803), .C(n56), .Z(n2155) );
  COND1XL U2609 ( .A(n2767), .B(n1861), .C(n2127), .Z(n878) );
  CANR2X1 U2610 ( .A(result[41]), .B(n2758), .C(n2752), .D(n2662), .Z(n2127)
         );
  COND1XL U2611 ( .A(n2767), .B(n1860), .C(n2131), .Z(n874) );
  CANR2X1 U2612 ( .A(result[45]), .B(n2758), .C(n2752), .D(n2665), .Z(n2131)
         );
  COND1XL U2613 ( .A(n2767), .B(n2676), .C(n2129), .Z(n876) );
  CANR2X1 U2614 ( .A(result[43]), .B(n2758), .C(n2752), .D(n2666), .Z(n2129)
         );
  COND1XL U2615 ( .A(n2767), .B(n1858), .C(n2135), .Z(n870) );
  CANR2X1 U2616 ( .A(result[49]), .B(n2758), .C(n2752), .D(n2674), .Z(n2135)
         );
  COND1XL U2617 ( .A(n2768), .B(n1857), .C(n2137), .Z(n868) );
  CANR2X1 U2618 ( .A(result[51]), .B(n2758), .C(n2752), .D(n2675), .Z(n2137)
         );
  COND1XL U2619 ( .A(n2767), .B(n2679), .C(n2133), .Z(n872) );
  CANR2X1 U2620 ( .A(result[47]), .B(n2758), .C(n2752), .D(n2670), .Z(n2133)
         );
  COND1XL U2621 ( .A(n112), .B(n2768), .C(n2139), .Z(n866) );
  CANR2X1 U2622 ( .A(result[53]), .B(n2757), .C(n2751), .D(n2678), .Z(n2139)
         );
  CANR2X1 U2623 ( .A(result[55]), .B(n2757), .C(n2751), .D(n2681), .Z(n2141)
         );
  COND1XL U2624 ( .A(n108), .B(n2769), .C(n2143), .Z(n862) );
  CANR2X1 U2625 ( .A(result[57]), .B(n2757), .C(n2751), .D(n2682), .Z(n2143)
         );
  CANR2X1 U2626 ( .A(result[59]), .B(n2757), .C(n2751), .D(n2683), .Z(n2145)
         );
  COND1XL U2627 ( .A(n104), .B(n2769), .C(n2147), .Z(n858) );
  CANR2X1 U2628 ( .A(result[61]), .B(n2757), .C(n2751), .D(n1984), .Z(n2147)
         );
  COND1XL U2629 ( .A(n102), .B(n2769), .C(n2647), .Z(n793) );
  CANR2X1 U2630 ( .A(result[63]), .B(n2757), .C(n2751), .D(n1851), .Z(n2647)
         );
  CND3XL U2631 ( .A(n53), .B(n1993), .C(n56), .Z(n1998) );
  CEOX1 U2632 ( .A(n2168), .B(n1982), .Z(n2164) );
  CANR5CXL U2633 ( .A(result[33]), .B(n2169), .C(n2156), .Z(n2168) );
  COND11X1 U2634 ( .A(n1994), .B(i[17]), .C(n2036), .D(n2037), .Z(n937) );
  CND2X1 U2635 ( .A(i[17]), .B(n2038), .Z(n2037) );
  COND11X1 U2636 ( .A(n2745), .B(i[21]), .C(n2046), .D(n2047), .Z(n933) );
  CND2X1 U2637 ( .A(i[21]), .B(n2048), .Z(n2047) );
  COND2X1 U2638 ( .A(n2003), .B(n1986), .C(n2745), .D(n2004), .Z(n951) );
  CND2X1 U2639 ( .A(i[0]), .B(n1986), .Z(n2004) );
  COND2X1 U2640 ( .A(n1985), .B(n2743), .C(i[0]), .D(n1994), .Z(n952) );
  COND1XL U2641 ( .A(n2763), .B(n1928), .C(n2091), .Z(n914) );
  CANR2X1 U2642 ( .A(result[5]), .B(n2761), .C(n2755), .D(n1838), .Z(n2091) );
  COND1XL U2643 ( .A(n2763), .B(n1921), .C(n2093), .Z(n912) );
  CANR2X1 U2644 ( .A(result[7]), .B(n2761), .C(n2755), .D(n1837), .Z(n2093) );
  COND1XL U2645 ( .A(n2764), .B(n1919), .C(n2099), .Z(n906) );
  CANR2X1 U2646 ( .A(result[13]), .B(n2761), .C(n2755), .D(n1848), .Z(n2099)
         );
  COND1XL U2647 ( .A(n2764), .B(n1918), .C(n2097), .Z(n908) );
  CANR2X1 U2648 ( .A(result[11]), .B(n2761), .C(n2755), .D(n1849), .Z(n2097)
         );
  COND1XL U2649 ( .A(n2763), .B(n2685), .C(n2095), .Z(n910) );
  CANR2X1 U2650 ( .A(result[9]), .B(n2761), .C(n2755), .D(n1850), .Z(n2095) );
  COND1XL U2651 ( .A(n2765), .B(n1909), .C(n2107), .Z(n898) );
  CANR2X1 U2652 ( .A(result[21]), .B(n2760), .C(n2754), .D(n1844), .Z(n2107)
         );
  COND1XL U2653 ( .A(n2764), .B(n1908), .C(n2105), .Z(n900) );
  CANR2X1 U2654 ( .A(result[19]), .B(n2760), .C(n2754), .D(n1845), .Z(n2105)
         );
  COND1XL U2655 ( .A(n2764), .B(n1906), .C(n2101), .Z(n904) );
  CANR2X1 U2656 ( .A(result[15]), .B(n2761), .C(n2755), .D(n1847), .Z(n2101)
         );
  COND1XL U2657 ( .A(n2764), .B(n1902), .C(n2103), .Z(n902) );
  CANR2X1 U2658 ( .A(result[17]), .B(n2760), .C(n2754), .D(n1846), .Z(n2103)
         );
  COND1XL U2659 ( .A(n2765), .B(n1896), .C(n2111), .Z(n894) );
  CANR2X1 U2660 ( .A(result[25]), .B(n2760), .C(n2754), .D(n1842), .Z(n2111)
         );
  COND1XL U2661 ( .A(n2765), .B(n1892), .C(n2113), .Z(n892) );
  CANR2X1 U2662 ( .A(result[27]), .B(n2760), .C(n2754), .D(n1841), .Z(n2113)
         );
  COND1XL U2663 ( .A(n2765), .B(n1888), .C(n2109), .Z(n896) );
  CANR2X1 U2664 ( .A(result[23]), .B(n2760), .C(n2754), .D(n1843), .Z(n2109)
         );
  COND1XL U2665 ( .A(n2765), .B(n1882), .C(n2115), .Z(n890) );
  CANR2X1 U2666 ( .A(result[29]), .B(n2759), .C(n2753), .D(n1836), .Z(n2115)
         );
  COND1XL U2667 ( .A(n2766), .B(n1881), .C(n2117), .Z(n888) );
  CANR2X1 U2668 ( .A(result[31]), .B(n2759), .C(n2753), .D(n2684), .Z(n2117)
         );
  COND1XL U2669 ( .A(n2766), .B(n2667), .C(n2119), .Z(n886) );
  COND1XL U2670 ( .A(n2766), .B(n1864), .C(n2121), .Z(n884) );
  CANR2X1 U2671 ( .A(result[35]), .B(n2759), .C(n2753), .D(n2660), .Z(n2121)
         );
  COND1XL U2672 ( .A(n2766), .B(n2671), .C(n2125), .Z(n880) );
  CANR2X1 U2673 ( .A(result[39]), .B(n2759), .C(n2753), .D(n2663), .Z(n2125)
         );
  COND1XL U2674 ( .A(n2766), .B(n1862), .C(n2123), .Z(n882) );
  CANR2X1 U2675 ( .A(result[37]), .B(n2759), .C(n2753), .D(n2661), .Z(n2123)
         );
  COND1XL U2676 ( .A(n2766), .B(n1967), .C(n2116), .Z(n889) );
  CANR2X1 U2677 ( .A(result[30]), .B(n2759), .C(n2753), .D(n1821), .Z(n2116)
         );
  COND1XL U2678 ( .A(n2766), .B(n1966), .C(n2118), .Z(n887) );
  COND1XL U2679 ( .A(n2763), .B(n1964), .C(n2090), .Z(n915) );
  CANR2X1 U2680 ( .A(result[4]), .B(n2761), .C(n2755), .D(n1833), .Z(n2090) );
  COND1XL U2681 ( .A(n2763), .B(n1963), .C(n2092), .Z(n913) );
  CANR2X1 U2682 ( .A(result[6]), .B(n2761), .C(n2755), .D(n1832), .Z(n2092) );
  COND1XL U2683 ( .A(n2763), .B(n1962), .C(n2094), .Z(n911) );
  CANR2X1 U2684 ( .A(result[8]), .B(n2761), .C(n2755), .D(n1835), .Z(n2094) );
  COND1XL U2685 ( .A(n2764), .B(n1961), .C(n2096), .Z(n909) );
  CANR2X1 U2686 ( .A(result[10]), .B(n2761), .C(n2755), .D(n1831), .Z(n2096)
         );
  COND1XL U2687 ( .A(n2764), .B(n1960), .C(n2098), .Z(n907) );
  CANR2X1 U2688 ( .A(result[12]), .B(n2761), .C(n2755), .D(n1830), .Z(n2098)
         );
  COND1XL U2689 ( .A(n2764), .B(n1959), .C(n2100), .Z(n905) );
  CANR2X1 U2690 ( .A(result[14]), .B(n2761), .C(n2755), .D(n1829), .Z(n2100)
         );
  COND1XL U2691 ( .A(n2764), .B(n1958), .C(n2102), .Z(n903) );
  CANR2X1 U2692 ( .A(result[16]), .B(n2760), .C(n2754), .D(n1828), .Z(n2102)
         );
  COND1XL U2693 ( .A(n2764), .B(n1957), .C(n2104), .Z(n901) );
  CANR2X1 U2694 ( .A(result[18]), .B(n2760), .C(n2754), .D(n1827), .Z(n2104)
         );
  COND1XL U2695 ( .A(n2765), .B(n1956), .C(n2106), .Z(n899) );
  CANR2X1 U2696 ( .A(result[20]), .B(n2760), .C(n2754), .D(n1826), .Z(n2106)
         );
  COND1XL U2697 ( .A(n2765), .B(n1955), .C(n2108), .Z(n897) );
  CANR2X1 U2698 ( .A(result[22]), .B(n2760), .C(n2754), .D(n1825), .Z(n2108)
         );
  COND1XL U2699 ( .A(n2765), .B(n1954), .C(n2110), .Z(n895) );
  CANR2X1 U2700 ( .A(result[24]), .B(n2760), .C(n2754), .D(n1824), .Z(n2110)
         );
  COND1XL U2701 ( .A(n2765), .B(n1953), .C(n2112), .Z(n893) );
  CANR2X1 U2702 ( .A(result[26]), .B(n2760), .C(n2754), .D(n1823), .Z(n2112)
         );
  COND1XL U2703 ( .A(n2765), .B(n1952), .C(n2114), .Z(n891) );
  CANR2X1 U2704 ( .A(result[28]), .B(n2759), .C(n2753), .D(n1822), .Z(n2114)
         );
  COND1XL U2705 ( .A(n2766), .B(n1951), .C(n2120), .Z(n885) );
  CANR2X1 U2706 ( .A(result[34]), .B(n2759), .C(n2753), .D(n1982), .Z(n2120)
         );
  COND1XL U2707 ( .A(n2766), .B(n1950), .C(n2122), .Z(n883) );
  CANR2X1 U2708 ( .A(result[36]), .B(n2759), .C(n2753), .D(n1981), .Z(n2122)
         );
  COND1XL U2709 ( .A(n2766), .B(n1949), .C(n2124), .Z(n881) );
  CANR2X1 U2710 ( .A(result[38]), .B(n2759), .C(n2753), .D(n1980), .Z(n2124)
         );
  COND1XL U2711 ( .A(n2767), .B(n1948), .C(n2126), .Z(n879) );
  CANR2X1 U2712 ( .A(result[40]), .B(n2758), .C(n2752), .D(n1979), .Z(n2126)
         );
  COND1XL U2713 ( .A(n2767), .B(n1947), .C(n2128), .Z(n877) );
  CANR2X1 U2714 ( .A(result[42]), .B(n2758), .C(n2752), .D(n1978), .Z(n2128)
         );
  COND1XL U2715 ( .A(n2767), .B(n1946), .C(n2130), .Z(n875) );
  CANR2X1 U2716 ( .A(result[44]), .B(n2758), .C(n2752), .D(n1977), .Z(n2130)
         );
  COND1XL U2717 ( .A(n2767), .B(n1945), .C(n2132), .Z(n873) );
  CANR2X1 U2718 ( .A(result[46]), .B(n2758), .C(n2752), .D(n1976), .Z(n2132)
         );
  COND1XL U2719 ( .A(n2767), .B(n1944), .C(n2134), .Z(n871) );
  CANR2X1 U2720 ( .A(result[48]), .B(n2758), .C(n2752), .D(n1975), .Z(n2134)
         );
  COND1XL U2721 ( .A(n2768), .B(n1943), .C(n2136), .Z(n869) );
  CANR2X1 U2722 ( .A(result[50]), .B(n2758), .C(n2752), .D(n1974), .Z(n2136)
         );
  COND1XL U2723 ( .A(n2768), .B(n1942), .C(n2138), .Z(n867) );
  CANR2X1 U2724 ( .A(result[52]), .B(n2757), .C(n2751), .D(n1973), .Z(n2138)
         );
  COND1XL U2725 ( .A(n2768), .B(n1941), .C(n2140), .Z(n865) );
  CANR2X1 U2726 ( .A(result[54]), .B(n2757), .C(n2751), .D(n1972), .Z(n2140)
         );
  COND1XL U2727 ( .A(n2768), .B(n1940), .C(n2142), .Z(n863) );
  CANR2X1 U2728 ( .A(result[56]), .B(n2757), .C(n2751), .D(n1971), .Z(n2142)
         );
  COND1XL U2729 ( .A(n2768), .B(n1939), .C(n2144), .Z(n861) );
  CANR2X1 U2730 ( .A(result[58]), .B(n2757), .C(n2751), .D(n1970), .Z(n2144)
         );
  COND1XL U2731 ( .A(n2768), .B(n1938), .C(n2146), .Z(n859) );
  CANR2X1 U2732 ( .A(result[60]), .B(n2757), .C(n2751), .D(n1969), .Z(n2146)
         );
  COND1XL U2733 ( .A(n2768), .B(n1937), .C(n2148), .Z(n857) );
  CANR2X1 U2734 ( .A(result[62]), .B(n2757), .C(n2751), .D(n1983), .Z(n2148)
         );
  COND1XL U2735 ( .A(n1802), .B(n2686), .C(n1987), .Z(n957) );
  CANR2X1 U2736 ( .A(n1988), .B(n1989), .C(nst[0]), .D(n1799), .Z(n1987) );
  COND4CX1 U2737 ( .A(n2003), .B(n2005), .C(n1930), .D(n2006), .Z(n950) );
  CND4X1 U2738 ( .A(n2771), .B(i[1]), .C(i[0]), .D(n1930), .Z(n2006) );
  CND2X1 U2739 ( .A(n2770), .B(n1986), .Z(n2005) );
  COND4CX1 U2740 ( .A(n2000), .B(n2009), .C(n1924), .D(n2010), .Z(n948) );
  CND4X1 U2741 ( .A(n2771), .B(i[5]), .C(n2002), .D(n1924), .Z(n2010) );
  CND2X1 U2742 ( .A(n2770), .B(n1926), .Z(n2009) );
  COND4CX1 U2743 ( .A(n1996), .B(n2007), .C(n1923), .D(n2008), .Z(n949) );
  CND4X1 U2744 ( .A(n2771), .B(i[3]), .C(n1999), .D(n1923), .Z(n2008) );
  CND2X1 U2745 ( .A(n2770), .B(n1925), .Z(n2007) );
  COND4CX1 U2746 ( .A(n2011), .B(n2014), .C(n1915), .D(n2015), .Z(n946) );
  CND4X1 U2747 ( .A(n2771), .B(i[7]), .C(n2013), .D(n1915), .Z(n2015) );
  CND2X1 U2748 ( .A(n2770), .B(n1917), .Z(n2014) );
  COND4CX1 U2749 ( .A(n2016), .B(n2019), .C(n1914), .D(n2020), .Z(n944) );
  CND4X1 U2750 ( .A(n2771), .B(i[9]), .C(n2018), .D(n1914), .Z(n2020) );
  CND2X1 U2751 ( .A(n2770), .B(n1916), .Z(n2019) );
  COND4CX1 U2752 ( .A(n2026), .B(n2029), .C(n1900), .D(n2030), .Z(n940) );
  CND4X1 U2753 ( .A(n2771), .B(i[13]), .C(n2028), .D(n1900), .Z(n2030) );
  CND2X1 U2754 ( .A(n2770), .B(n1901), .Z(n2029) );
  COND4CX1 U2755 ( .A(n2021), .B(n2024), .C(n1897), .D(n2025), .Z(n942) );
  CND4X1 U2756 ( .A(n2771), .B(i[11]), .C(n2023), .D(n1897), .Z(n2025) );
  CND2X1 U2757 ( .A(n2770), .B(n1920), .Z(n2024) );
  COND4CX1 U2758 ( .A(n2031), .B(n2033), .C(n1895), .D(n2034), .Z(n938) );
  CND2X1 U2759 ( .A(n2770), .B(n1899), .Z(n2033) );
  COND4CX1 U2760 ( .A(n2041), .B(n2043), .C(n1874), .D(n2044), .Z(n934) );
  CND2X1 U2761 ( .A(n2771), .B(n1893), .Z(n2043) );
  CND2X1 U2762 ( .A(n2039), .B(n2040), .Z(n936) );
  CND4X1 U2763 ( .A(n2771), .B(i[17]), .C(n1894), .D(n1885), .Z(n2040) );
  COND4CX1 U2764 ( .A(n2770), .B(n1886), .C(n2038), .D(i[18]), .Z(n2039) );
  CND2X1 U2765 ( .A(n2049), .B(n2050), .Z(n932) );
  COND4CX1 U2766 ( .A(n2770), .B(n1879), .C(n2048), .D(i[22]), .Z(n2049) );
  CENX1 U2767 ( .A(opera1[30]), .B(n2782), .Z(n2353) );
  CND2X1 U2768 ( .A(valid), .B(n1988), .Z(n2076) );
  CND2X1 U2769 ( .A(n1990), .B(n1797), .Z(n1992) );
  CNR2X1 U2770 ( .A(n2707), .B(nst[0]), .Z(n55) );
  CEOXL U2771 ( .A(n2334), .B(n2335), .Z(n2329) );
  CEOXL U2772 ( .A(n2346), .B(n2347), .Z(n2345) );
  CEOXL U2773 ( .A(n2270), .B(n2271), .Z(n2269) );
  CEOXL U2774 ( .A(n2245), .B(n2246), .Z(n2244) );
  CEOXL U2775 ( .A(n2320), .B(n2321), .Z(n2319) );
  CEOXL U2776 ( .A(n2295), .B(n2296), .Z(n2294) );
  CEOXL U2777 ( .A(n2194), .B(n2195), .Z(n2193) );
  CEOXL U2778 ( .A(opera1[29]), .B(n2777), .Z(n2446) );
  CEOXL U2779 ( .A(opera1[28]), .B(n2777), .Z(n2444) );
  CEOX1 U2780 ( .A(n2166), .B(n2167), .Z(n2389) );
  CND3XL U2781 ( .A(n2394), .B(n2167), .C(n2166), .Z(n2395) );
  COND4CXL U2782 ( .A(res_not_wire[22]), .B(n1903), .C(n987), .D(n2592), .Z(
        n2586) );
  COND4CXL U2783 ( .A(res_not_wire[12]), .B(n1912), .C(n978), .D(n2532), .Z(
        n2526) );
  COND4CXL U2784 ( .A(res_not_wire[16]), .B(n1907), .C(n984), .D(n2556), .Z(
        n2550) );
  COND4CXL U2785 ( .A(res_not_wire[14]), .B(n1911), .C(n983), .D(n2544), .Z(
        n2538) );
  COND4CXL U2786 ( .A(res_not_wire[60]), .B(n2333), .C(n1852), .D(n2086), .Z(
        n2341) );
  COND4CXL U2787 ( .A(res_not_wire[44]), .B(n2233), .C(n995), .D(n2247), .Z(
        n2241) );
  COND4CXL U2788 ( .A(res_not_wire[48]), .B(n2258), .C(n997), .D(n2272), .Z(
        n2266) );
  CEOXL U2789 ( .A(res_not_wire[14]), .B(n2532), .Z(n2533) );
  CEOXL U2790 ( .A(res_not_wire[18]), .B(n2556), .Z(n2557) );
  CEOXL U2791 ( .A(n2333), .B(n1938), .Z(n2336) );
  CEOXL U2792 ( .A(n2233), .B(n1946), .Z(n2236) );
  CEOXL U2793 ( .A(n2258), .B(n1944), .Z(n2261) );
  CANR4CXL U2794 ( .A(n2322), .B(n1939), .C(n106), .D(n2333), .Z(n2332) );
  CANR4CXL U2795 ( .A(n2222), .B(n1947), .C(n2676), .D(n2233), .Z(n2232) );
  CANR4CXL U2796 ( .A(n2247), .B(n1945), .C(n2679), .D(n2258), .Z(n2257) );
  COND4CXL U2797 ( .A(res_not_wire[24]), .B(n1891), .C(n985), .D(n2604), .Z(
        n2598) );
  COND4CXL U2798 ( .A(res_not_wire[20]), .B(n1904), .C(n981), .D(n2580), .Z(
        n2574) );
  COND4CXL U2799 ( .A(res_not_wire[2]), .B(n1934), .C(n975), .D(n2472), .Z(
        n2466) );
  COND4CXL U2800 ( .A(res_not_wire[6]), .B(n2489), .C(n977), .D(n2496), .Z(
        n2490) );
  COND4CXL U2801 ( .A(res_not_wire[56]), .B(n2308), .C(n1853), .D(n2322), .Z(
        n2316) );
  COND4CXL U2802 ( .A(res_not_wire[52]), .B(n2283), .C(n1855), .D(n2297), .Z(
        n2291) );
  COND4CXL U2803 ( .A(res_not_wire[40]), .B(n2207), .C(n994), .D(n2222), .Z(
        n2216) );
  COND4CXL U2804 ( .A(res_not_wire[36]), .B(n2181), .C(n993), .D(n2196), .Z(
        n2190) );
  CEOXL U2805 ( .A(res_not_wire[26]), .B(n2604), .Z(n2605) );
  CEOXL U2806 ( .A(res_not_wire[22]), .B(n2580), .Z(n2581) );
  CEOXL U2807 ( .A(n2472), .B(n2701), .Z(n2473) );
  CEOXL U2808 ( .A(n2308), .B(n1940), .Z(n2311) );
  CEOXL U2809 ( .A(n2283), .B(n1942), .Z(n2286) );
  CEOXL U2810 ( .A(n2207), .B(n1948), .Z(n2210) );
  CEOXL U2811 ( .A(n2181), .B(n1950), .Z(n2184) );
  CANR4CXL U2812 ( .A(n2297), .B(n1941), .C(n110), .D(n2308), .Z(n2307) );
  CANR4CXL U2813 ( .A(n2272), .B(n1943), .C(n1857), .D(n2283), .Z(n2282) );
  CANR4CXL U2814 ( .A(n2196), .B(n1949), .C(n2671), .D(n2207), .Z(n2206) );
  CANR4CXL U2815 ( .A(n1870), .B(n1951), .C(n1864), .D(n2181), .Z(n2180) );
  CIVX1 U2816 ( .A(n2655), .Z(n2750) );
  CIVXL U2817 ( .A(n2657), .Z(n2769) );
  CIVXL U2818 ( .A(n2784), .Z(n2778) );
  CIVXL U2819 ( .A(n2784), .Z(n2779) );
  CIVXL U2820 ( .A(n2784), .Z(n2780) );
  CIVXL U2821 ( .A(n2783), .Z(n2781) );
  CIVXL U2822 ( .A(n2784), .Z(n2782) );
endmodule


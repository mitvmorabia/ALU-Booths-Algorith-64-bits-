
module multiplier ( result, valid, opera1, opera2, muordi, clock, reset, start
 );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input muordi, clock, reset, start;
  output valid;
  wire   opera2_63, N34, n18, n38, n43, n52, n53, n55, n56, n108, n114, n116,
         n118, n120, n122, n126, n128, n130, n132, n134, n136, n138, n142,
         n144, n146, n148, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n1125, n1126, n1128, n1138, n1472, n1473, n1474, n1475,
         n1476, n1849, n1891, n1918, n2060, n2276, n2281, n2284, n2298, n2309,
         n2313, n2314, n2315, n2316, n2321, n2322, n2323, n2324, n2327, n2329,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2343, n2345,
         n2346, n2347, n2348, n2350, n2351, n2352, n2353, n2354, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2372, n2379, n2380, n2382, n2391, n2393, n2396, n2397,
         n2408, n2418, n2424, n2435, n2439, n2531, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2570, n2574, n2576,
         n2581, n2583, n2585, n2588, n2590, n2591, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n3153, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661;
  wire   [63:0] res_not_wire;
  wire   [2:0] nst;
  wire   [31:0] i;
  tri   c_inop1;
  tri   c_inop2;
  tri   c_inres;
  assign opera2_63 = opera2[63];

  CTSX2 A3 ( .A(1'b1), .E(n3511), .Z(c_inop2) );
  CTSX2 A2 ( .A(1'b0), .E(n3313), .Z(c_inop1) );
  CFD1QX2 \i_reg[26]  ( .D(n3267), .CP(clock), .Q(i[26]) );
  CFD2X1 \cst_reg[2]  ( .D(N34), .CP(clock), .CD(n2276), .Q(n3433), .QN(n2060)
         );
  CIVX2 U1724 ( .A(i[29]), .Z(n2281) );
  CIVX2 U1727 ( .A(i[26]), .Z(n2284) );
  CIVX2 U1741 ( .A(i[10]), .Z(n2298) );
  CIVX2 U1756 ( .A(res_not_wire[44]), .Z(n2313) );
  CIVX2 U1757 ( .A(res_not_wire[56]), .Z(n2314) );
  CIVX2 U1758 ( .A(res_not_wire[8]), .Z(n2315) );
  CIVX2 U1759 ( .A(res_not_wire[58]), .Z(n2316) );
  CIVX2 U1764 ( .A(n1128), .Z(n2321) );
  CIVX2 U1765 ( .A(n1126), .Z(n2322) );
  CIVX2 U1766 ( .A(n1125), .Z(n2323) );
  CIVX2 U1767 ( .A(n3396), .Z(n2324) );
  CIVX2 U1770 ( .A(result[51]), .Z(n2327) );
  CIVX2 U1779 ( .A(nst[2]), .Z(n2336) );
  CIVX2 U1780 ( .A(nst[1]), .Z(n2337) );
  CIVX2 U1782 ( .A(result[19]), .Z(n2339) );
  CIVX2 U1783 ( .A(result[30]), .Z(n2340) );
  CIVX2 U1784 ( .A(result[29]), .Z(n2341) );
  CIVX2 U1786 ( .A(result[21]), .Z(n2343) );
  CIVX2 U1788 ( .A(result[15]), .Z(n2345) );
  CIVX2 U1789 ( .A(result[23]), .Z(n2346) );
  CIVX2 U1791 ( .A(result[7]), .Z(n2348) );
  CIVX2 U1793 ( .A(result[9]), .Z(n2350) );
  CIVX2 U1794 ( .A(result[5]), .Z(n2351) );
  CIVX2 U1795 ( .A(result[3]), .Z(n2352) );
  CIVX2 U1796 ( .A(result[1]), .Z(n2353) );
  CIVX2 U1797 ( .A(result[22]), .Z(n2354) );
  CIVX2 U1799 ( .A(result[28]), .Z(n2356) );
  CIVX2 U1800 ( .A(result[24]), .Z(n2357) );
  CIVX2 U1801 ( .A(result[16]), .Z(n2358) );
  CIVX2 U1802 ( .A(result[12]), .Z(n2359) );
  CIVX2 U1803 ( .A(result[10]), .Z(n2360) );
  CIVX2 U1804 ( .A(result[6]), .Z(n2361) );
  CIVX2 U1805 ( .A(result[4]), .Z(n2362) );
  CIVX2 U1806 ( .A(result[2]), .Z(n2363) );
  CIVX2 U1807 ( .A(result[11]), .Z(n2364) );
  CIVX2 U1808 ( .A(result[14]), .Z(n2365) );
  CIVX2 U1809 ( .A(result[8]), .Z(n2366) );
  CIVX2 U1810 ( .A(result[26]), .Z(n2367) );
  CIVX2 U1811 ( .A(result[20]), .Z(n2368) );
  CIVX2 U1815 ( .A(res_not_wire[62]), .Z(n2372) );
  CIVX2 U1822 ( .A(result[57]), .Z(n2379) );
  CIVX2 U1825 ( .A(n1473), .Z(n2382) );
  CIVX2 U1839 ( .A(res_not_wire[10]), .Z(n2396) );
  CIVX2 U1840 ( .A(res_not_wire[14]), .Z(n2397) );
  CIVX2 U1861 ( .A(result[53]), .Z(n2418) );
  CIVX2 U1867 ( .A(res_not_wire[30]), .Z(n2424) );
  CND2IX1 U1934 ( .B(n3288), .A(nst[1]), .Z(n52) );
  CTSX2 A1 ( .A(1'b1), .E(opera1[31]), .Z(c_inop1) );
  CFD1QXL \result_reg[55]  ( .D(n833), .CP(clock), .Q(result[55]) );
  CFD1QXL \result_reg[51]  ( .D(n837), .CP(clock), .Q(result[51]) );
  CFD1QXL \result_reg[57]  ( .D(n831), .CP(clock), .Q(result[57]) );
  CFD1QXL \nst_reg[2]  ( .D(n921), .CP(clock), .Q(nst[2]) );
  CFD1QXL \nst_reg[1]  ( .D(n922), .CP(clock), .Q(nst[1]) );
  CFD1QXL \nst_reg[0]  ( .D(n3161), .CP(clock), .Q(nst[0]) );
  CFD1QXL \res_not_reg[63]  ( .D(n793), .CP(clock), .Q(n1476) );
  CFD1QXL \result_reg[24]  ( .D(n801), .CP(clock), .Q(result[24]) );
  CFD1XL \res_not_reg[62]  ( .D(n857), .CP(clock), .Q(res_not_wire[62]), .QN(
        n3223) );
  CFD1QXL \result_reg[19]  ( .D(n3270), .CP(clock), .Q(result[19]) );
  CFD1QXL \result_reg[30]  ( .D(n795), .CP(clock), .Q(result[30]) );
  CFD1QXL \result_reg[29]  ( .D(n796), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[27]  ( .D(n798), .CP(clock), .Q(result[27]) );
  CFD1QXL \result_reg[21]  ( .D(n804), .CP(clock), .Q(result[21]) );
  CFD1QXL \result_reg[17]  ( .D(n808), .CP(clock), .Q(result[17]) );
  CFD1QXL \result_reg[15]  ( .D(n3274), .CP(clock), .Q(result[15]) );
  CFD1QXL \result_reg[23]  ( .D(n802), .CP(clock), .Q(result[23]) );
  CFD1QXL \result_reg[7]  ( .D(n3162), .CP(clock), .Q(result[7]) );
  CFD1QXL \result_reg[13]  ( .D(n3275), .CP(clock), .Q(result[13]) );
  CFD1QXL \result_reg[9]  ( .D(n3276), .CP(clock), .Q(result[9]) );
  CFD1QXL \result_reg[5]  ( .D(n3261), .CP(clock), .Q(result[5]) );
  CFD1QXL \result_reg[1]  ( .D(n3277), .CP(clock), .Q(result[1]) );
  CFD1QXL \result_reg[22]  ( .D(n803), .CP(clock), .Q(result[22]) );
  CFD1QXL \result_reg[18]  ( .D(n807), .CP(clock), .Q(result[18]) );
  CFD1QXL \result_reg[28]  ( .D(n797), .CP(clock), .Q(result[28]) );
  CFD1QXL \result_reg[16]  ( .D(n809), .CP(clock), .Q(result[16]) );
  CFD1QXL \result_reg[12]  ( .D(n3279), .CP(clock), .Q(result[12]) );
  CFD1QXL \result_reg[10]  ( .D(n3163), .CP(clock), .Q(result[10]) );
  CFD1QXL \result_reg[6]  ( .D(n3280), .CP(clock), .Q(result[6]) );
  CFD1QXL \result_reg[2]  ( .D(n3281), .CP(clock), .Q(result[2]) );
  CFD1QXL \result_reg[11]  ( .D(n3282), .CP(clock), .Q(result[11]) );
  CFD1QXL \result_reg[14]  ( .D(n811), .CP(clock), .Q(result[14]) );
  CFD1QXL \result_reg[8]  ( .D(n3164), .CP(clock), .Q(result[8]) );
  CFD1QXL \result_reg[26]  ( .D(n799), .CP(clock), .Q(result[26]) );
  CFD1QXL \result_reg[20]  ( .D(n805), .CP(clock), .Q(result[20]) );
  CFD1QXL \result_reg[3]  ( .D(n3283), .CP(clock), .Q(result[3]) );
  CFD1XL \res_not_reg[61]  ( .D(n858), .CP(clock), .Q(n1126), .QN(n3251) );
  CFD1QXL \result_reg[4]  ( .D(n821), .CP(clock), .Q(result[4]) );
  CFD1QXL \result_reg[63]  ( .D(n919), .CP(clock), .Q(result[63]) );
  CFD1XL \res_not_reg[30]  ( .D(n889), .CP(clock), .Q(res_not_wire[30]), .QN(
        n3190) );
  CFD1XL \res_not_reg[54]  ( .D(n865), .CP(clock), .Q(res_not_wire[54]) );
  CFD1XL \res_not_reg[59]  ( .D(n860), .CP(clock), .Q(n1125), .QN(n3222) );
  CFD1XL \res_not_reg[58]  ( .D(n861), .CP(clock), .Q(res_not_wire[58]), .QN(
        n3250) );
  CFD1QXL \result_reg[0]  ( .D(n3284), .CP(clock), .Q(result[0]) );
  CFD1QXL \res_not_reg[26]  ( .D(n893), .CP(clock), .Q(res_not_wire[26]) );
  CFD1XL \res_not_reg[48]  ( .D(n871), .CP(clock), .Q(res_not_wire[48]) );
  CFD1QXL \res_not_reg[9]  ( .D(n910), .CP(clock), .Q(n1474) );
  CFD1XL \res_not_reg[24]  ( .D(n895), .CP(clock), .Q(res_not_wire[24]), .QN(
        n3176) );
  CFD1XL \res_not_reg[44]  ( .D(n875), .CP(clock), .Q(res_not_wire[44]), .QN(
        n3187) );
  CFD1XL \res_not_reg[53]  ( .D(n866), .CP(clock), .Q(n1128) );
  CFD1QXL \i_reg[31]  ( .D(n955), .CP(clock), .Q(i[31]) );
  CFD1XL \res_not_reg[45]  ( .D(n874), .CP(clock), .Q(n3236), .QN(n120) );
  CFD1XL \res_not_reg[29]  ( .D(n890), .CP(clock), .QN(n136) );
  CFD1XL \res_not_reg[12]  ( .D(n907), .CP(clock), .Q(res_not_wire[12]), .QN(
        n3378) );
  CFD1QXL \res_not_reg[11]  ( .D(n908), .CP(clock), .Q(n1918) );
  CFD1XL \res_not_reg[27]  ( .D(n892), .CP(clock), .QN(n138) );
  CFD1XL \res_not_reg[17]  ( .D(n902), .CP(clock), .QN(n148) );
  CFD1XL \res_not_reg[43]  ( .D(n876), .CP(clock), .Q(n3220), .QN(n122) );
  CFD1XL \res_not_reg[49]  ( .D(n870), .CP(clock), .Q(n3226), .QN(n116) );
  CTSX2 A5 ( .A(1'b1), .E(n18), .Z(c_inres) );
  CTSX2 A6 ( .A(1'b0), .E(n3541), .Z(c_inres) );
  CFD1XL \res_not_reg[14]  ( .D(n905), .CP(clock), .Q(res_not_wire[14]), .QN(
        n3247) );
  CFD1XL \res_not_reg[8]  ( .D(n911), .CP(clock), .Q(res_not_wire[8]), .QN(
        n3248) );
  CFD1XL \res_not_reg[18]  ( .D(n901), .CP(clock), .Q(res_not_wire[18]), .QN(
        n3188) );
  CFD1XL \res_not_reg[28]  ( .D(n891), .CP(clock), .Q(res_not_wire[28]) );
  CFD1XL \res_not_reg[15]  ( .D(n904), .CP(clock), .Q(n43), .QN(n3189) );
  CFD1X1 \res_not_reg[2]  ( .D(n917), .CP(clock), .Q(res_not_wire[2]) );
  CFD1QXL \res_not_reg[7]  ( .D(n912), .CP(clock), .Q(n1891) );
  CFD1X1 \res_not_reg[0]  ( .D(n920), .CP(clock), .Q(res_not_wire[0]) );
  CFD1X1 \res_not_reg[20]  ( .D(n899), .CP(clock), .Q(res_not_wire[20]) );
  CFD1XL \res_not_reg[46]  ( .D(n873), .CP(clock), .Q(res_not_wire[46]), .QN(
        n3237) );
  CFD1QXL \res_not_reg[13]  ( .D(n906), .CP(clock), .Q(n1475) );
  CFD1XL \res_not_reg[10]  ( .D(n909), .CP(clock), .Q(res_not_wire[10]), .QN(
        n3253) );
  CFD1XL \res_not_reg[50]  ( .D(n869), .CP(clock), .Q(res_not_wire[50]), .QN(
        n3256) );
  CFD1XL \res_not_reg[52]  ( .D(n867), .CP(clock), .Q(res_not_wire[52]), .QN(
        n3257) );
  CFD1QX1 \i_reg[22]  ( .D(n932), .CP(clock), .Q(i[22]) );
  CFD1XL \result_reg[41]  ( .D(n847), .CP(clock), .Q(result[41]), .QN(n3184)
         );
  CFD1XL \result_reg[35]  ( .D(n853), .CP(clock), .Q(result[35]), .QN(n3439)
         );
  CFD1XL \result_reg[50]  ( .D(n838), .CP(clock), .Q(result[50]), .QN(n3299)
         );
  CFD1XL \result_reg[38]  ( .D(n850), .CP(clock), .Q(result[38]), .QN(n3424)
         );
  CFD1XL \res_not_reg[40]  ( .D(n879), .CP(clock), .Q(res_not_wire[40]), .QN(
        n3255) );
  CFD1XL \result_reg[52]  ( .D(n836), .CP(clock), .Q(result[52]), .QN(n3311)
         );
  CFD1XL \res_not_reg[16]  ( .D(n903), .CP(clock), .Q(res_not_wire[16]), .QN(
        n3241) );
  CFD1XL \result_reg[34]  ( .D(n854), .CP(clock), .Q(result[34]), .QN(n3178)
         );
  CFD1XL \result_reg[44]  ( .D(n844), .CP(clock), .Q(result[44]), .QN(n3221)
         );
  CFD1XL \result_reg[36]  ( .D(n852), .CP(clock), .Q(result[36]) );
  CFD1XL \result_reg[39]  ( .D(n849), .CP(clock), .Q(result[39]), .QN(n3249)
         );
  CFD1XL \result_reg[43]  ( .D(n845), .CP(clock), .Q(result[43]), .QN(n3244)
         );
  CFD1XL \result_reg[40]  ( .D(n848), .CP(clock), .Q(result[40]) );
  CFD1XL \result_reg[37]  ( .D(n851), .CP(clock), .Q(result[37]), .QN(n3442)
         );
  CFD1X1 \result_reg[46]  ( .D(n842), .CP(clock), .Q(result[46]) );
  CFD1XL \res_not_reg[51]  ( .D(n868), .CP(clock), .QN(n114) );
  CFD1XL \res_not_reg[60]  ( .D(n859), .CP(clock), .Q(res_not_wire[60]), .QN(
        n3171) );
  CFD1QX1 \result_reg[47]  ( .D(n841), .CP(clock), .Q(result[47]) );
  CFD1XL \res_not_reg[41]  ( .D(n878), .CP(clock), .Q(n3234), .QN(n3185) );
  CFD1X1 \res_not_reg[6]  ( .D(n913), .CP(clock), .Q(res_not_wire[6]), .QN(
        n3183) );
  CFD1QXL \result_reg[32]  ( .D(n856), .CP(clock), .Q(result[32]) );
  CFD1XL \result_reg[42]  ( .D(n846), .CP(clock), .Q(result[42]) );
  CFD1QX1 \result_reg[31]  ( .D(n794), .CP(clock), .Q(result[31]) );
  CFD1XL \result_reg[48]  ( .D(n840), .CP(clock), .Q(result[48]), .QN(n3321)
         );
  CFD1XL \res_not_reg[23]  ( .D(n896), .CP(clock), .QN(n142) );
  CFD1XL \res_not_reg[39]  ( .D(n880), .CP(clock), .Q(n3173), .QN(n126) );
  CFD1XL \res_not_reg[21]  ( .D(n898), .CP(clock), .QN(n144) );
  CFD1XL \res_not_reg[37]  ( .D(n882), .CP(clock), .Q(n3174), .QN(n128) );
  CFD1XL \res_not_reg[57]  ( .D(n862), .CP(clock), .QN(n108) );
  CFD1XL \res_not_reg[56]  ( .D(n863), .CP(clock), .Q(res_not_wire[56]), .QN(
        n3224) );
  CFD1XL \res_not_reg[55]  ( .D(n864), .CP(clock), .Q(n1138), .QN(n3252) );
  CFD1XL \res_not_reg[25]  ( .D(n894), .CP(clock), .Q(n38), .QN(n3229) );
  CFD1XL \res_not_reg[35]  ( .D(n884), .CP(clock), .QN(n130) );
  CFD1XL \res_not_reg[42]  ( .D(n877), .CP(clock), .Q(res_not_wire[42]) );
  CFD1QXL \i_reg[5]  ( .D(n953), .CP(clock), .Q(i[5]) );
  CFD1XL \res_not_reg[22]  ( .D(n897), .CP(clock), .Q(res_not_wire[22]), .QN(
        n3180) );
  CFD1QX1 \result_reg[25]  ( .D(n800), .CP(clock), .Q(result[25]) );
  CFD1QX1 \result_reg[61]  ( .D(n827), .CP(clock), .Q(result[61]) );
  CFD1QX1 \result_reg[54]  ( .D(n834), .CP(clock), .Q(result[54]) );
  CFD1QX1 \result_reg[53]  ( .D(n835), .CP(clock), .Q(result[53]) );
  CFD1QX1 \i_reg[28]  ( .D(n926), .CP(clock), .Q(i[28]) );
  CFD1QX1 \i_reg[11]  ( .D(n943), .CP(clock), .Q(i[11]) );
  CFD1QX1 \i_reg[25]  ( .D(n929), .CP(clock), .Q(i[25]) );
  CFD1QX1 \i_reg[24]  ( .D(n930), .CP(clock), .Q(i[24]) );
  CFD4X1 \cst_reg[0]  ( .D(n55), .CP(clock), .SD(n2276), .Q(n56), .QN(n3513)
         );
  CFD1XL \res_not_reg[31]  ( .D(n888), .CP(clock), .Q(n3789), .QN(n134) );
  CFD1QXL valid_reg ( .D(n923), .CP(clock), .Q(valid) );
  CFD1X1 sign_reg ( .D(n3290), .CP(clock), .Q(n18), .QN(n3541) );
  CFD1QX1 \res_not_reg[5]  ( .D(n914), .CP(clock), .Q(n1473) );
  CFD1QX1 \i_reg[18]  ( .D(n936), .CP(clock), .Q(i[18]) );
  CFD1QX1 \result_reg[62]  ( .D(n826), .CP(clock), .Q(result[62]) );
  CFD1XL \res_not_reg[38]  ( .D(n881), .CP(clock), .Q(res_not_wire[38]), .QN(
        n3258) );
  CFD1XL \res_not_reg[47]  ( .D(n872), .CP(clock), .Q(n3254), .QN(n118) );
  CFD1XL \result_reg[33]  ( .D(n855), .CP(clock), .Q(result[33]), .QN(n3242)
         );
  CFD1XL \res_not_reg[36]  ( .D(n883), .CP(clock), .Q(res_not_wire[36]), .QN(
        n3240) );
  CFD1XL \res_not_reg[19]  ( .D(n900), .CP(clock), .Q(n3230), .QN(n146) );
  CFD1X1 \res_not_reg[4]  ( .D(n915), .CP(clock), .Q(res_not_wire[4]), .QN(
        n3225) );
  CFD1QX1 \i_reg[30]  ( .D(n3168), .CP(clock), .Q(i[30]) );
  CFD1QX1 \i_reg[27]  ( .D(n927), .CP(clock), .Q(i[27]) );
  CFD1QX1 \i_reg[23]  ( .D(n931), .CP(clock), .Q(i[23]) );
  CFD1QX1 \i_reg[20]  ( .D(n934), .CP(clock), .Q(i[20]) );
  CFD1QX1 \i_reg[19]  ( .D(n935), .CP(clock), .Q(i[19]) );
  CFD1QX1 \i_reg[15]  ( .D(n939), .CP(clock), .Q(i[15]) );
  CFD1QX1 \i_reg[12]  ( .D(n942), .CP(clock), .Q(i[12]) );
  CFD1QX1 \i_reg[10]  ( .D(n944), .CP(clock), .Q(i[10]) );
  CFD1QX1 \i_reg[9]  ( .D(n945), .CP(clock), .Q(i[9]) );
  CFD1QX1 \i_reg[7]  ( .D(n947), .CP(clock), .Q(i[7]) );
  CFD1QX1 \i_reg[6]  ( .D(n948), .CP(clock), .Q(i[6]) );
  CFD1QX1 \i_reg[2]  ( .D(n950), .CP(clock), .Q(i[2]) );
  CFD1QX1 \i_reg[1]  ( .D(n951), .CP(clock), .Q(i[1]) );
  CFD1QX1 \i_reg[0]  ( .D(n3265), .CP(clock), .Q(i[0]) );
  CFD1QX1 \res_not_reg[3]  ( .D(n916), .CP(clock), .Q(n1472) );
  CFD1QX1 \i_reg[3]  ( .D(n3262), .CP(clock), .Q(i[3]) );
  CFD1QXL \i_reg[4]  ( .D(n949), .CP(clock), .Q(i[4]) );
  CFD1QX1 \res_not_reg[1]  ( .D(n918), .CP(clock), .Q(n1849) );
  CFD1QX1 \res_not_reg[34]  ( .D(n885), .CP(clock), .Q(n3396) );
  CFD1XL \i_reg[8]  ( .D(n946), .CP(clock), .Q(n3373), .QN(n3374) );
  CFD1QXL \res_not_reg[32]  ( .D(n887), .CP(clock), .Q(n3349) );
  CFD1QX1 \result_reg[56]  ( .D(n832), .CP(clock), .Q(result[56]) );
  CTSX2 A4 ( .A(1'b0), .E(n3194), .Z(c_inop2) );
  CFD1QXL \i_reg[16]  ( .D(n938), .CP(clock), .Q(i[16]) );
  CFD1QX1 \result_reg[60]  ( .D(n4659), .CP(clock), .Q(result[60]) );
  CFD1QX1 \result_reg[45]  ( .D(n843), .CP(clock), .Q(result[45]) );
  CFD1XL \res_not_reg[33]  ( .D(n3263), .CP(clock), .Q(n3198), .QN(n132) );
  CFD1QX1 \i_reg[21]  ( .D(n933), .CP(clock), .Q(i[21]) );
  CFD1QX1 \i_reg[17]  ( .D(n3169), .CP(clock), .Q(i[17]) );
  CFD1QX1 \i_reg[14]  ( .D(n940), .CP(clock), .Q(i[14]) );
  CFD1QX1 \i_reg[13]  ( .D(n941), .CP(clock), .Q(i[13]) );
  CFD1X1 \result_reg[49]  ( .D(n839), .CP(clock), .Q(result[49]), .QN(n3177)
         );
  CFD1QX2 \result_reg[59]  ( .D(n829), .CP(clock), .Q(result[59]) );
  CFD4XL \cst_reg[1]  ( .D(n52), .CP(clock), .SD(n2276), .Q(n53), .QN(n3545)
         );
  CFD1QX1 \i_reg[29]  ( .D(n3268), .CP(clock), .Q(i[29]) );
  CFD1QX1 \result_reg[58]  ( .D(n830), .CP(clock), .Q(result[58]) );
  CNIVX1 U1935 ( .A(n957), .Z(n3161) );
  CNIVX1 U1936 ( .A(n818), .Z(n3162) );
  CND2IX2 U1937 ( .B(n3406), .A(n4249), .Z(n4250) );
  CENXL U1938 ( .A(opera2[27]), .B(n3197), .Z(n4344) );
  CND3X1 U1939 ( .A(n4375), .B(n4272), .C(n4190), .Z(n4196) );
  CNIVX1 U1940 ( .A(n815), .Z(n3163) );
  CNIVX1 U1941 ( .A(n817), .Z(n3164) );
  CNIVXL U1942 ( .A(n4120), .Z(n3165) );
  CENX1 U1943 ( .A(n3440), .B(n4245), .Z(n4169) );
  CNIVX1 U1944 ( .A(n4169), .Z(n3166) );
  COND1X2 U1945 ( .A(n3509), .B(n2393), .C(n2531), .Z(n920) );
  CIVXL U1946 ( .A(res_not_wire[20]), .Z(n2435) );
  CMXI2X2 U1947 ( .A0(n4630), .A1(n4629), .S(i[25]), .Z(n929) );
  CNIVX1 U1948 ( .A(result[47]), .Z(n3167) );
  CNIVX1 U1949 ( .A(n924), .Z(n3168) );
  CMXI2XL U1950 ( .A0(n4651), .A1(n4650), .S(i[30]), .Z(n924) );
  CMX2XL U1951 ( .A0(n4608), .A1(n4611), .S(i[20]), .Z(n934) );
  CMXI2X2 U1952 ( .A0(n4578), .A1(n4577), .S(i[10]), .Z(n944) );
  CMXI2X2 U1953 ( .A0(n4574), .A1(n4573), .S(i[9]), .Z(n945) );
  CMXI2X2 U1954 ( .A0(n4562), .A1(n3445), .S(i[2]), .Z(n950) );
  CMXI2X2 U1955 ( .A0(n4561), .A1(n3453), .S(i[1]), .Z(n951) );
  CMXI2X2 U1956 ( .A0(n4614), .A1(n4613), .S(i[21]), .Z(n933) );
  CNIVX1 U1957 ( .A(n937), .Z(n3169) );
  CMXI2X2 U1958 ( .A0(n4592), .A1(n4591), .S(i[13]), .Z(n941) );
  CEOX4 U1959 ( .A(opera1[0]), .B(opera1[31]), .Z(n3444) );
  CANR1X1 U1960 ( .A(n3983), .B(n4400), .C(n3989), .Z(n3984) );
  CND3X2 U1961 ( .A(n4288), .B(n4287), .C(n4286), .Z(n4362) );
  CANR1X2 U1962 ( .A(n3652), .B(n3651), .C(n3337), .Z(n3343) );
  CND2X1 U1963 ( .A(n3434), .B(n4505), .Z(n3332) );
  CIVDX4 U1964 ( .A(opera2_63), .Z0(n3196), .Z1(n3197) );
  CNR2XL U1965 ( .A(n4067), .B(n4066), .Z(n4068) );
  CND2X2 U1966 ( .A(n4502), .B(n3305), .Z(n3809) );
  CND2X2 U1967 ( .A(n3213), .B(result[51]), .Z(n4502) );
  CND2X2 U1968 ( .A(n3192), .B(n4488), .Z(n3836) );
  CND2X2 U1969 ( .A(n4545), .B(n3835), .Z(n3775) );
  CAN2X2 U1970 ( .A(n3655), .B(n3690), .Z(n3300) );
  CND2X2 U1971 ( .A(n3477), .B(n3444), .Z(n3663) );
  CEOX2 U1972 ( .A(opera1[18]), .B(opera1[31]), .Z(n3415) );
  CND2X1 U1973 ( .A(n3838), .B(n3338), .Z(n3804) );
  CIVX1 U1974 ( .A(n3809), .Z(n3491) );
  CND2X2 U1975 ( .A(n3300), .B(result[48]), .Z(n3835) );
  CEOX4 U1976 ( .A(opera1[9]), .B(opera1[31]), .Z(n3486) );
  CNR2IXL U1977 ( .B(n3352), .A(n3358), .Z(n3699) );
  COAN1X1 U1978 ( .A(n3352), .B(n3709), .C(n3708), .Z(n3323) );
  CND2XL U1979 ( .A(n3684), .B(n3676), .Z(n3677) );
  CNR2X2 U1980 ( .A(n3682), .B(n3684), .Z(n3615) );
  CNIVX4 U1981 ( .A(opera1[31]), .Z(n3215) );
  CND2X2 U1982 ( .A(n3614), .B(n3451), .Z(n3683) );
  CNR2IXL U1983 ( .B(n3451), .A(n3682), .Z(n3667) );
  CND2XL U1984 ( .A(n3669), .B(n3670), .Z(n3671) );
  CNR3X1 U1985 ( .A(n3990), .B(n3989), .C(n4028), .Z(n3991) );
  COND1X1 U1986 ( .A(n4553), .B(n4416), .C(n4415), .Z(n830) );
  CEOX4 U1987 ( .A(opera1[15]), .B(n3353), .Z(n3688) );
  CIVX20 U1988 ( .A(opera1[31]), .Z(n3353) );
  CND2X1 U1989 ( .A(n4410), .B(n4397), .Z(n3982) );
  CND2X1 U1990 ( .A(n3848), .B(n3849), .Z(n3653) );
  CANR1X1 U1991 ( .A(n4402), .B(n4065), .C(n3982), .Z(n3989) );
  CND2X1 U1992 ( .A(n3611), .B(n3548), .Z(n3514) );
  CND2IX1 U1993 ( .B(n3980), .A(n3383), .Z(n3384) );
  CENX2 U1994 ( .A(opera1[3]), .B(opera1[31]), .Z(n3555) );
  CND3X1 U1995 ( .A(n3615), .B(n3616), .C(n3617), .Z(n3631) );
  CNR2X1 U1996 ( .A(n3673), .B(n3631), .Z(n3621) );
  CEOX2 U1997 ( .A(opera1[10]), .B(opera1[31]), .Z(n3352) );
  COAN1X1 U1998 ( .A(n3414), .B(n3306), .C(n3651), .Z(n3213) );
  CNR2IX1 U1999 ( .B(n4042), .A(n4044), .Z(n3403) );
  CEOX2 U2000 ( .A(opera1[2]), .B(opera1[31]), .Z(n3477) );
  CND2X1 U2001 ( .A(n3298), .B(n3805), .Z(n3964) );
  CND2IX1 U2002 ( .B(n3311), .A(n3343), .Z(n3848) );
  CND2X1 U2003 ( .A(n3213), .B(result[51]), .Z(n3475) );
  CND4X1 U2004 ( .A(c_inres), .B(n3218), .C(n4176), .D(res_not_wire[6]), .Z(
        n4278) );
  CNIVX2 U2005 ( .A(opera2_63), .Z(n3195) );
  CND4X1 U2006 ( .A(n4161), .B(n4097), .C(n4096), .D(n4095), .Z(n4261) );
  CND2X1 U2007 ( .A(n3993), .B(n3992), .Z(n3995) );
  CND2X1 U2008 ( .A(n3335), .B(n3336), .Z(n4383) );
  CNIVX1 U2009 ( .A(n4457), .Z(n3340) );
  CND2X1 U2010 ( .A(c_inop2), .B(n4080), .Z(n4234) );
  CND3XL U2011 ( .A(n1891), .B(res_not_wire[8]), .C(n3588), .Z(n4262) );
  CND2X1 U2012 ( .A(res_not_wire[24]), .B(n4122), .Z(n4380) );
  CANR1X1 U2013 ( .A(n4420), .B(n3813), .C(n3812), .Z(n3814) );
  CENX1 U2014 ( .A(n1138), .B(n4422), .Z(n3818) );
  CENX1 U2015 ( .A(result[63]), .B(n4034), .Z(n4039) );
  CND2X1 U2016 ( .A(n3384), .B(n3385), .Z(n4416) );
  CND2IX4 U2017 ( .B(n3358), .A(n3317), .Z(n3711) );
  COAN1X1 U2018 ( .A(n3437), .B(n3756), .C(n3755), .Z(n3758) );
  CND2IX1 U2019 ( .B(n3748), .A(result[60]), .Z(n4053) );
  CND2IX1 U2020 ( .B(n4345), .A(n4208), .Z(n4353) );
  CNR3X1 U2021 ( .A(n114), .B(n3852), .C(n3968), .Z(n3879) );
  CAN2X1 U2022 ( .A(n3436), .B(n3433), .Z(n4394) );
  CAN3X2 U2023 ( .A(n3435), .B(n3635), .C(n3427), .Z(n3754) );
  COND4CX1 U2024 ( .A(n3213), .B(result[51]), .C(n3765), .D(n3434), .Z(n3806)
         );
  CNR2X1 U2025 ( .A(n3513), .B(n3433), .Z(n3432) );
  CND2IX2 U2026 ( .B(n3752), .A(result[59]), .Z(n3985) );
  CEOX1 U2027 ( .A(result[61]), .B(n3744), .Z(n4052) );
  CENX1 U2028 ( .A(opera2[4]), .B(opera2_63), .Z(n3170) );
  CIVX2 U2029 ( .A(n3170), .Z(n3440) );
  CND4X1 U2030 ( .A(n3597), .B(n4089), .C(n3596), .D(n3595), .Z(n4363) );
  CNR4X1 U2031 ( .A(i[1]), .B(i[2]), .C(i[3]), .D(i[0]), .Z(n3532) );
  CND2IX1 U2032 ( .B(n4381), .A(n4382), .Z(n3336) );
  CENX1 U2033 ( .A(n3204), .B(n4546), .Z(n4554) );
  CND2XL U2034 ( .A(n3634), .B(n3621), .Z(n3655) );
  CAN2X1 U2035 ( .A(n3927), .B(n3867), .Z(n4476) );
  CND2X1 U2036 ( .A(n3980), .B(n3985), .Z(n3482) );
  COR2X1 U2037 ( .A(n3970), .B(n116), .Z(n3852) );
  CND2IX1 U2038 ( .B(n3171), .A(n4046), .Z(n4045) );
  CEOX1 U2039 ( .A(opera2[6]), .B(opera2_63), .Z(n3199) );
  CND6X2 U2040 ( .A(n1918), .B(res_not_wire[10]), .C(n1474), .D(n1891), .E(
        res_not_wire[8]), .F(n3588), .Z(n4191) );
  CND2IX1 U2041 ( .B(n4327), .A(n3233), .Z(n4372) );
  CNR5XL U2042 ( .A(n3237), .B(n118), .C(n4365), .D(n134), .E(n4480), .Z(n3408) );
  CND2XL U2043 ( .A(n3433), .B(n3545), .Z(n3546) );
  CND2IX1 U2044 ( .B(n4384), .A(n4383), .Z(n4388) );
  CND2IX1 U2045 ( .B(n3664), .A(n3665), .Z(n3658) );
  CENX1 U2046 ( .A(n3747), .B(n3628), .Z(n3744) );
  CENX1 U2047 ( .A(result[59]), .B(n3752), .Z(n3172) );
  CIVX2 U2048 ( .A(n3172), .Z(n3980) );
  CAN4X1 U2049 ( .A(res_not_wire[38]), .B(res_not_wire[42]), .C(n3173), .D(
        n3174), .Z(n3422) );
  CEOX1 U2050 ( .A(opera2[5]), .B(opera2_63), .Z(n3328) );
  CND4X1 U2051 ( .A(n4090), .B(n4123), .C(res_not_wire[18]), .D(
        res_not_wire[16]), .Z(n4209) );
  COAN1X1 U2052 ( .A(n4645), .B(i[1]), .C(n3453), .Z(n3445) );
  CND4X1 U2053 ( .A(n4571), .B(n4582), .C(i[12]), .D(i[13]), .Z(n4594) );
  CEOX1 U2054 ( .A(result[54]), .B(n3764), .Z(n3846) );
  CND2IX1 U2055 ( .B(n4382), .A(n4381), .Z(n3335) );
  CND2X1 U2056 ( .A(result[33]), .B(n3401), .Z(n3922) );
  CMXI2XL U2057 ( .A0(n4652), .A1(n3413), .S(result[60]), .Z(n2597) );
  CEOX1 U2058 ( .A(result[39]), .B(n3722), .Z(n3942) );
  CND2X1 U2059 ( .A(n3242), .B(n3915), .Z(n3567) );
  CAN3X2 U2060 ( .A(n3410), .B(n4024), .C(n4023), .Z(n4031) );
  CNR2XL U2061 ( .A(n4027), .B(n3763), .Z(n3781) );
  CNR3XL U2062 ( .A(n128), .B(n3941), .C(n126), .Z(n3412) );
  COND3X1 U2063 ( .A(n3964), .B(n3809), .C(n3807), .D(n3808), .Z(n3847) );
  CNR2X1 U2064 ( .A(n3250), .B(n3222), .Z(n3421) );
  CAN4X1 U2065 ( .A(i[18]), .B(i[19]), .C(i[22]), .D(i[23]), .Z(n3575) );
  CNR4X1 U2066 ( .A(n3852), .B(n4365), .C(n3851), .D(n3853), .Z(n4537) );
  CND4X1 U2067 ( .A(n4118), .B(n4112), .C(n4114), .D(n4113), .Z(n4345) );
  CND2IX1 U2068 ( .B(n4326), .A(res_not_wire[18]), .Z(n4370) );
  CNR2IX1 U2069 ( .B(result[47]), .A(n4495), .Z(n4497) );
  CMXI2XL U2070 ( .A0(n4652), .A1(n3413), .S(result[13]), .Z(n2550) );
  CEOX1 U2071 ( .A(opera1[8]), .B(opera1[31]), .Z(n3479) );
  CND3X1 U2072 ( .A(n3622), .B(n3634), .C(n3621), .Z(n3657) );
  CND2XL U2073 ( .A(n3677), .B(n3687), .Z(n3678) );
  CND2X1 U2074 ( .A(n3184), .B(n3723), .Z(n3726) );
  CAOR1X1 U2075 ( .A(n3558), .B(n3557), .C(n3368), .Z(n3175) );
  CIVX2 U2076 ( .A(n3175), .Z(n3228) );
  CNR2X1 U2077 ( .A(n3176), .B(n3180), .Z(n3591) );
  CND2X1 U2078 ( .A(n3373), .B(i[9]), .Z(n4575) );
  CANR2XL U2079 ( .A(n3410), .B(n4024), .C(n3629), .D(result[61]), .Z(n3316)
         );
  CANR11X1 U2080 ( .A(n4477), .B(n3867), .C(n3927), .D(n3689), .Z(n3838) );
  CND4X1 U2081 ( .A(i[25]), .B(i[26]), .C(i[14]), .D(i[27]), .Z(n3578) );
  CND2XL U2082 ( .A(res_not_wire[12]), .B(n4089), .Z(n4269) );
  CNR2XL U2083 ( .A(n3513), .B(n3545), .Z(n3436) );
  CNR2XL U2084 ( .A(n3497), .B(n4046), .Z(n3999) );
  CNR2IX1 U2085 ( .B(i[20]), .A(n4609), .Z(n3456) );
  CANR1X1 U2086 ( .A(n3216), .B(n3878), .C(n3346), .Z(n3850) );
  CND2X2 U2087 ( .A(n4291), .B(n3789), .Z(n3968) );
  CIVX2 U2088 ( .A(n4365), .Z(n4291) );
  COR2X1 U2089 ( .A(n4280), .B(n4175), .Z(n4135) );
  COR2X1 U2090 ( .A(n4115), .B(n4338), .Z(n4226) );
  CND2IXL U2091 ( .B(n4625), .A(i[16]), .Z(n4599) );
  COND3XL U2092 ( .A(n3863), .B(n4466), .C(n3864), .D(n3862), .Z(n3902) );
  CMXI2XL U2093 ( .A0(n4652), .A1(n3413), .S(result[18]), .Z(n2555) );
  CIVXL U2094 ( .A(n3644), .Z(n3306) );
  COR2X1 U2095 ( .A(n3723), .B(n3184), .Z(n3725) );
  CND2IX2 U2096 ( .B(n3706), .A(result[55]), .Z(n4042) );
  CND2X1 U2097 ( .A(n4475), .B(n3679), .Z(n3680) );
  CAN3X2 U2098 ( .A(n3705), .B(n4476), .C(n3899), .Z(n3297) );
  COR2X1 U2099 ( .A(n3774), .B(n3177), .Z(n4545) );
  CND4X1 U2100 ( .A(res_not_wire[44]), .B(n3871), .C(n3220), .D(n3236), .Z(
        n4480) );
  CND2X1 U2101 ( .A(result[36]), .B(n3228), .Z(n3733) );
  CND2X1 U2102 ( .A(n3178), .B(n3570), .Z(n4442) );
  CNR2IX1 U2103 ( .B(n3440), .A(n4245), .Z(n3406) );
  CNR2X1 U2104 ( .A(n3252), .B(n3224), .Z(n3243) );
  CND4X1 U2105 ( .A(n3373), .B(i[9]), .C(i[10]), .D(i[11]), .Z(n4588) );
  CND4X1 U2106 ( .A(n4631), .B(n4632), .C(i[25]), .D(i[24]), .Z(n4640) );
  CANR1XL U2107 ( .A(n4294), .B(n3500), .C(n3401), .Z(n4295) );
  CENX1 U2108 ( .A(result[53]), .B(n3777), .Z(n3216) );
  CNR2X1 U2109 ( .A(n4151), .B(n4152), .Z(n4101) );
  COR2X1 U2110 ( .A(n4318), .B(n3189), .Z(n4324) );
  CNR3XL U2111 ( .A(n3180), .B(n4222), .C(n142), .Z(n3202) );
  CND2IX1 U2112 ( .B(n4363), .A(res_not_wire[30]), .Z(n4365) );
  CND2IXL U2113 ( .B(n4625), .A(n3456), .Z(n4614) );
  CENX1 U2116 ( .A(n4514), .B(n126), .Z(n4527) );
  CMXI2XL U2117 ( .A0(n4652), .A1(n3413), .S(result[27]), .Z(n2564) );
  CNR2IX1 U2118 ( .B(n3480), .A(n4052), .Z(n3410) );
  CND2X1 U2119 ( .A(n4520), .B(n4519), .Z(n3825) );
  COND3X1 U2120 ( .A(n3179), .B(n3802), .C(n3860), .D(n3862), .Z(n3833) );
  CIVX2 U2121 ( .A(n3803), .Z(n3179) );
  COND1X1 U2122 ( .A(n3300), .B(result[48]), .C(n3835), .Z(n4487) );
  CND3X1 U2123 ( .A(result[46]), .B(n3677), .C(n3687), .Z(n4475) );
  CND2XL U2124 ( .A(n3221), .B(n3693), .Z(n3694) );
  CND2X1 U2125 ( .A(n3439), .B(n3569), .Z(n4440) );
  COR4X1 U2126 ( .A(n3433), .B(n2276), .C(n3545), .D(n3513), .Z(n3548) );
  CIVXL U2127 ( .A(reset), .Z(n2276) );
  COND1X1 U2128 ( .A(n4504), .B(n4503), .C(n3475), .Z(n4505) );
  CNR2X1 U2129 ( .A(n3224), .B(n108), .Z(n3231) );
  CNR2X1 U2130 ( .A(n4399), .B(n4043), .Z(n4051) );
  CIVX2 U2131 ( .A(n3777), .Z(n3649) );
  COND1XL U2132 ( .A(n116), .B(n3972), .C(n3256), .Z(n3973) );
  CND3XL U2133 ( .A(n3199), .B(n3328), .C(n3406), .Z(n4175) );
  CND2X1 U2134 ( .A(n3378), .B(n4191), .Z(n4192) );
  CNR2X1 U2135 ( .A(n3180), .B(n4302), .Z(n4305) );
  CND3X1 U2136 ( .A(n4118), .B(n4117), .C(n4116), .Z(n4338) );
  CIVX2 U2137 ( .A(n4374), .Z(n4118) );
  COR2X1 U2138 ( .A(n4586), .B(n3374), .Z(n4574) );
  CNR2XL U2139 ( .A(n4609), .B(n4625), .Z(n4608) );
  COR2X1 U2140 ( .A(n4647), .B(n2281), .Z(n4651) );
  CND3XL U2141 ( .A(n4394), .B(n4495), .C(n4514), .Z(n3953) );
  CMXI2X1 U2142 ( .A0(n4652), .A1(n3413), .S(result[17]), .Z(n2554) );
  CND3XL U2143 ( .A(n3181), .B(n4345), .C(n4121), .Z(n4129) );
  CIVX2 U2144 ( .A(n4384), .Z(n3181) );
  CND2IX1 U2145 ( .B(n3663), .A(n3666), .Z(n3673) );
  CND4X1 U2146 ( .A(n3675), .B(n3659), .C(n3686), .D(n3685), .Z(n3768) );
  CAN8X1 U2147 ( .A(n3635), .B(n3488), .C(n3437), .D(n3435), .E(n3429), .F(
        n3428), .G(n3427), .H(n3182), .Z(n3238) );
  CIVXL U2148 ( .A(n3630), .Z(n3182) );
  CND2IX1 U2149 ( .B(n3747), .A(n3627), .Z(n4015) );
  CND2IX1 U2150 ( .B(result[45]), .A(n3681), .Z(n3867) );
  CND4X1 U2151 ( .A(n1474), .B(n1891), .C(res_not_wire[8]), .D(n3588), .Z(
        n4264) );
  CNR2XL U2152 ( .A(n3990), .B(n3989), .Z(n3986) );
  COR2X1 U2153 ( .A(n3480), .B(n4421), .Z(n3474) );
  CEOX1 U2154 ( .A(n3915), .B(n3242), .Z(n3916) );
  CND2X1 U2155 ( .A(n118), .B(n4494), .Z(n4498) );
  CENX1 U2156 ( .A(n3424), .B(n3446), .Z(n3423) );
  CANR2X1 U2157 ( .A(result[39]), .B(n3721), .C(n4517), .D(n4516), .Z(n4522)
         );
  COND3XL U2158 ( .A(n4446), .B(n4448), .C(n4445), .D(n4444), .Z(n4450) );
  COAN1X1 U2159 ( .A(n3301), .B(n3967), .C(n3305), .Z(n4504) );
  CAOR1X1 U2160 ( .A(res_not_wire[40]), .B(n3399), .C(n3234), .Z(n4455) );
  CND4X1 U2161 ( .A(res_not_wire[62]), .B(n1126), .C(res_not_wire[60]), .D(
        n4046), .Z(n4074) );
  COR4X1 U2162 ( .A(n4241), .B(n4242), .C(n4234), .D(n4233), .Z(n4245) );
  CND2IX1 U2163 ( .B(n4152), .A(n4099), .Z(n4189) );
  CND2X1 U2164 ( .A(n3183), .B(n4254), .Z(n4177) );
  CND3XL U2165 ( .A(n3309), .B(n4104), .C(n4145), .Z(n4317) );
  COR4X1 U2166 ( .A(n148), .B(n3241), .C(n3189), .D(n4318), .Z(n4326) );
  CND2XL U2167 ( .A(n3190), .B(n4363), .Z(n4364) );
  CND4XL U2168 ( .A(n3548), .B(n3547), .C(n3546), .D(n3583), .Z(n4391) );
  COND4CX1 U2169 ( .A(n4534), .B(n3243), .C(n108), .D(n3365), .Z(n4010) );
  CNR2XL U2170 ( .A(n4588), .B(n4586), .Z(n4583) );
  CNR2X1 U2171 ( .A(n4624), .B(n4625), .Z(n4621) );
  COND4CXL U2172 ( .A(res_not_wire[52]), .B(n3879), .C(n1128), .D(n3854), .Z(
        n3857) );
  CEOXL U2173 ( .A(res_not_wire[22]), .B(n4302), .Z(n4230) );
  CENX1 U2174 ( .A(opera1[14]), .B(opera1[31]), .Z(n3684) );
  CND3XL U2175 ( .A(n3667), .B(n3659), .C(n3675), .Z(n3669) );
  CND2X1 U2176 ( .A(n3317), .B(n3699), .Z(n3708) );
  CNR2XL U2177 ( .A(n3747), .B(n3628), .Z(n3354) );
  COAN1X1 U2178 ( .A(n3479), .B(n3715), .C(n3714), .Z(n3716) );
  CND2XL U2179 ( .A(n3184), .B(n3723), .Z(n3724) );
  CNR2X1 U2180 ( .A(n3255), .B(n3185), .Z(n3450) );
  CND3XL U2181 ( .A(n3186), .B(res_not_wire[2]), .C(n1849), .Z(n4167) );
  CIVX2 U2182 ( .A(n4231), .Z(n3186) );
  CND4X1 U2183 ( .A(n4105), .B(n3309), .C(n4104), .D(n4145), .Z(n4327) );
  CND2IX1 U2184 ( .B(n3653), .A(n3847), .Z(n4530) );
  COND3XL U2185 ( .A(n3925), .B(n3926), .C(n3680), .D(n3924), .Z(n3345) );
  CND4X1 U2186 ( .A(n4060), .B(n4057), .C(n4058), .D(n4059), .Z(n4067) );
  CND3XL U2187 ( .A(n4631), .B(i[21]), .C(n3456), .Z(n4616) );
  CND2X1 U2188 ( .A(n3240), .B(n4430), .Z(n3602) );
  COND1XL U2189 ( .A(n122), .B(n4469), .C(n3187), .Z(n3872) );
  COR3X2 U2190 ( .A(n3941), .B(n128), .C(n3968), .Z(n4514) );
  CENX1 U2191 ( .A(n4432), .B(n4431), .Z(n4433) );
  CND2XL U2192 ( .A(n3188), .B(n4326), .Z(n4218) );
  CEOXL U2193 ( .A(n4175), .B(n4280), .Z(n4281) );
  CND2XL U2194 ( .A(n3189), .B(n4318), .Z(n4319) );
  CNR2X1 U2195 ( .A(n3592), .B(n4370), .Z(n3404) );
  CND2IX1 U2196 ( .B(n3434), .A(n3331), .Z(n3333) );
  CND2IX1 U2197 ( .B(n4625), .A(n4626), .Z(n4630) );
  CND2IX1 U2198 ( .B(n4578), .A(i[10]), .Z(n4581) );
  CENX1 U2199 ( .A(n3846), .B(n3850), .Z(n3858) );
  CND2X1 U2200 ( .A(n3610), .B(n3227), .Z(n3607) );
  COND3XL U2201 ( .A(n3191), .B(n3840), .C(n3502), .D(n4544), .Z(n3845) );
  CIVX2 U2202 ( .A(n3839), .Z(n3191) );
  CMXI2XL U2203 ( .A0(n4652), .A1(n3413), .S(result[61]), .Z(n2598) );
  CENX1 U2204 ( .A(n4333), .B(n144), .Z(n4342) );
  CNR2XL U2205 ( .A(n2379), .B(n4495), .Z(n4009) );
  CIVX2 U2206 ( .A(n3722), .Z(n3721) );
  CIVX2 U2207 ( .A(n4487), .Z(n3192) );
  CIVXL U2208 ( .A(n4487), .Z(n4493) );
  CEOX1 U2209 ( .A(opera2[1]), .B(n3194), .Z(n4233) );
  CIVX16 U2210 ( .A(opera1[31]), .Z(n3296) );
  CIVX2 U2211 ( .A(n3695), .Z(n3659) );
  CIVX2 U2212 ( .A(n3483), .Z(n3987) );
  CENX2 U2213 ( .A(opera2[0]), .B(opera2_63), .Z(n4081) );
  CND2X4 U2214 ( .A(n3351), .B(n3470), .Z(n3664) );
  CENX4 U2215 ( .A(opera1[6]), .B(n3296), .Z(n3470) );
  CENXL U2216 ( .A(n3441), .B(n3944), .Z(n3582) );
  CIVXL U2217 ( .A(res_not_wire[4]), .Z(n2408) );
  CND4X2 U2218 ( .A(n3841), .B(n3792), .C(n3791), .D(res_not_wire[54]), .Z(
        n3815) );
  CND2IXL U2219 ( .B(n3237), .A(n3400), .Z(n4494) );
  CEOXL U2220 ( .A(res_not_wire[46]), .B(n3400), .Z(n3425) );
  CIVDX2 U2221 ( .A(opera2_63), .Z0(n3194), .Z1(n3193) );
  CIVX1 U2222 ( .A(n4422), .Z(n4534) );
  CIVX2 U2223 ( .A(n3353), .Z(n3512) );
  CIVX20 U2224 ( .A(opera1[31]), .Z(n3313) );
  CND3X2 U2225 ( .A(n4291), .B(n3793), .C(n3231), .Z(n4411) );
  CNR2IX2 U2226 ( .B(n1138), .A(n3815), .Z(n3793) );
  CENX1 U2227 ( .A(result[60]), .B(n3748), .Z(n3370) );
  CND2X1 U2228 ( .A(n3862), .B(n4466), .Z(n3705) );
  CND2X1 U2229 ( .A(result[60]), .B(n3200), .Z(n4057) );
  CENX1 U2230 ( .A(opera2[3]), .B(opera2_63), .Z(n4241) );
  CANR1XL U2231 ( .A(n4065), .B(n4064), .C(n4063), .Z(n4066) );
  CND2X1 U2232 ( .A(n3718), .B(n3293), .Z(n3696) );
  CIVX2 U2233 ( .A(n3658), .Z(n3660) );
  CIVX2 U2234 ( .A(n3664), .Z(n3718) );
  CENX1 U2235 ( .A(opera1[30]), .B(opera1[31]), .Z(n4013) );
  CIVX2 U2236 ( .A(n3703), .Z(n3704) );
  CND2X1 U2237 ( .A(n3834), .B(n3297), .Z(n3298) );
  CND2X1 U2238 ( .A(n3747), .B(n3746), .Z(n3748) );
  CND2X1 U2239 ( .A(result[43]), .B(n3704), .Z(n3862) );
  CND2X1 U2240 ( .A(result[39]), .B(n3721), .Z(n4515) );
  CNR2X1 U2241 ( .A(n3599), .B(n3598), .Z(n3585) );
  CNR2IX1 U2242 ( .B(n3417), .A(n4130), .Z(n4096) );
  CENX1 U2243 ( .A(opera2[7]), .B(n3197), .Z(n4280) );
  CND3X1 U2244 ( .A(n3591), .B(n3590), .C(n3589), .Z(n3592) );
  COND1XL U2245 ( .A(n3926), .B(n3925), .C(n3924), .Z(n3302) );
  CND2X1 U2246 ( .A(n4534), .B(n3243), .Z(n4425) );
  CENX1 U2247 ( .A(res_not_wire[58]), .B(n4411), .Z(n4414) );
  CNIVXL U2248 ( .A(n4503), .Z(n3322) );
  CENX1 U2249 ( .A(res_not_wire[4]), .B(n4252), .Z(n4168) );
  CENX1 U2250 ( .A(n4118), .B(n4336), .Z(n4107) );
  CENX1 U2251 ( .A(n4161), .B(n4242), .Z(n4162) );
  CND2X1 U2252 ( .A(n4101), .B(n4100), .Z(n4272) );
  CND2X1 U2253 ( .A(n4094), .B(n4093), .Z(n4243) );
  COND1XL U2254 ( .A(n4501), .B(n4553), .C(n4500), .Z(n841) );
  CANR4CX1 U2255 ( .A(n3334), .B(n4484), .C(n4483), .D(n4482), .Z(n4485) );
  CANR1XL U2256 ( .A(n3334), .B(n4484), .C(n4553), .Z(n4483) );
  CENX1 U2257 ( .A(n3216), .B(n3878), .Z(n3884) );
  CENX1 U2258 ( .A(n4286), .B(n4288), .Z(n4214) );
  CMX2X1 U2259 ( .A0(n3419), .A1(n4596), .S(i[14]), .Z(n940) );
  CMXI2XL U2260 ( .A0(n4599), .A1(n3454), .S(i[17]), .Z(n937) );
  CAN3X2 U2261 ( .A(n3510), .B(n4653), .C(n3541), .Z(n3413) );
  CIVX2 U2262 ( .A(n4495), .Z(n3200) );
  CAN2X1 U2263 ( .A(n4054), .B(n4065), .Z(n3201) );
  CIVX2 U2264 ( .A(n4553), .Z(n3502) );
  CIVXL U2265 ( .A(n1849), .Z(n3203) );
  CIVDX1 U2266 ( .A(n3497), .Z0(n3207), .Z1(n3208) );
  CIVDX1 U2267 ( .A(n3395), .Z0(n3211), .Z1(n3212) );
  CIVX2 U2268 ( .A(n3217), .Z(n3510) );
  CIVX1 U2269 ( .A(n3217), .Z(n3509) );
  COAN1X1 U2270 ( .A(result[52]), .B(n3766), .C(n3848), .Z(n3434) );
  CND3X1 U2271 ( .A(n1473), .B(res_not_wire[4]), .C(res_not_wire[0]), .Z(n3587) );
  CIVXL U2272 ( .A(n4547), .Z(n3204) );
  CIVX2 U2273 ( .A(n3204), .Z(n3205) );
  CIVX2 U2274 ( .A(n3773), .Z(n4547) );
  COND4CXL U2275 ( .A(n3837), .B(n3838), .C(n3836), .D(n3835), .Z(n3840) );
  CENX1 U2276 ( .A(opera2[8]), .B(opera2_63), .Z(n4134) );
  CND2XL U2277 ( .A(n3561), .B(n3444), .Z(n3565) );
  CIVX1 U2278 ( .A(n3771), .Z(n3643) );
  CND2IXL U2279 ( .B(result[50]), .A(n3771), .Z(n3772) );
  CNR3X1 U2280 ( .A(n3684), .B(n3683), .C(n3682), .Z(n3674) );
  CANR3X1 U2281 ( .A(n4051), .B(n4050), .C(n4048), .D(n4049), .Z(n4069) );
  CND2IX1 U2282 ( .B(n3839), .A(n3840), .Z(n4544) );
  CNR3X2 U2283 ( .A(n3375), .B(n3557), .C(n3555), .Z(n3206) );
  CNR3X2 U2284 ( .A(n3375), .B(n3557), .C(n3555), .Z(n3469) );
  CND2X2 U2285 ( .A(n3495), .B(n3238), .Z(n3755) );
  CIVX2 U2286 ( .A(n3196), .Z(n3511) );
  CND2XL U2287 ( .A(result[38]), .B(n3446), .Z(n3947) );
  CENX1 U2288 ( .A(n3424), .B(n3446), .Z(n3348) );
  CIVX1 U2289 ( .A(res_not_wire[22]), .Z(n2309) );
  CIVXL U2290 ( .A(n3349), .Z(n3350) );
  CND2X2 U2291 ( .A(c_inop1), .B(n3452), .Z(n3556) );
  COND1X1 U2292 ( .A(n3580), .B(n4594), .C(i[31]), .Z(n4512) );
  COND1X1 U2293 ( .A(n4553), .B(n4001), .C(n4000), .Z(n829) );
  CIVDXL U2294 ( .A(n3497), .Z0(n3209), .Z1(n3210) );
  CND3X1 U2295 ( .A(n3370), .B(n4007), .C(n3482), .Z(n4063) );
  CMXI2XL U2296 ( .A0(n3957), .A1(n3407), .S(i[4]), .Z(n949) );
  CMXI2XL U2297 ( .A0(n3610), .A1(n3607), .S(i[4]), .Z(n3608) );
  CNR2XL U2298 ( .A(i[19]), .B(i[4]), .Z(n3533) );
  CND2X1 U2299 ( .A(n4053), .B(n3201), .Z(n4047) );
  CND3X1 U2300 ( .A(n3584), .B(n4385), .C(n3583), .Z(n4495) );
  CND2X2 U2301 ( .A(opera1[7]), .B(n3313), .Z(n3356) );
  CIVX2 U2302 ( .A(n3688), .Z(n3617) );
  CND2X1 U2303 ( .A(n4515), .B(n3947), .Z(n3735) );
  CND2X1 U2304 ( .A(n3565), .B(n3564), .Z(n3915) );
  CND2X1 U2305 ( .A(res_not_wire[44]), .B(n3871), .Z(n3869) );
  CND2X1 U2306 ( .A(result[57]), .B(n3484), .Z(n4065) );
  CND3X1 U2307 ( .A(n3370), .B(n3759), .C(n3757), .Z(n4054) );
  CND2IX1 U2308 ( .B(n3392), .A(n4045), .Z(n4059) );
  COAN1X1 U2309 ( .A(n3471), .B(n3553), .C(n3730), .Z(n3446) );
  CND2X1 U2310 ( .A(n4515), .B(n3942), .Z(n4519) );
  CANR1X1 U2311 ( .A(n3304), .B(n3554), .C(n3553), .Z(n3728) );
  CND3X1 U2312 ( .A(res_not_wire[20]), .B(n3230), .C(n4334), .Z(n4222) );
  CIVX2 U2313 ( .A(n4353), .Z(n4288) );
  CND2X2 U2314 ( .A(n3584), .B(n3550), .Z(n4642) );
  CEOX2 U2315 ( .A(opera1[8]), .B(opera1[31]), .Z(n3493) );
  CENX1 U2316 ( .A(opera1[27]), .B(opera1[31]), .Z(n3749) );
  CENX1 U2317 ( .A(opera1[11]), .B(opera1[31]), .Z(n3682) );
  CND2X1 U2318 ( .A(n3559), .B(n3560), .Z(n3558) );
  CENX2 U2319 ( .A(opera1[31]), .B(opera1[4]), .Z(n3557) );
  CNR2X1 U2320 ( .A(i[21]), .B(i[20]), .Z(n3516) );
  CNR2X1 U2321 ( .A(i[24]), .B(i[23]), .Z(n3517) );
  CNR2X1 U2322 ( .A(i[10]), .B(i[9]), .Z(n3524) );
  CNR2X1 U2323 ( .A(i[7]), .B(i[6]), .Z(n3523) );
  CENX1 U2324 ( .A(opera1[28]), .B(opera1[31]), .Z(n3745) );
  CND2IX1 U2325 ( .B(n4474), .A(n3398), .Z(n3767) );
  COND1XL U2326 ( .A(n3560), .B(n3559), .C(n3558), .Z(n3569) );
  CND2X1 U2327 ( .A(n3428), .B(n3650), .Z(n3648) );
  CND2X1 U2328 ( .A(n3965), .B(n3772), .Z(n3773) );
  CND2X1 U2329 ( .A(n3396), .B(n4429), .Z(n3598) );
  CAOR1X1 U2330 ( .A(n3636), .B(n3638), .C(n3324), .Z(n3431) );
  CNR2IX1 U2331 ( .B(result[33]), .A(n3915), .Z(n3568) );
  CND3XL U2332 ( .A(i[14]), .B(i[15]), .C(n4593), .Z(n3552) );
  CND2IX1 U2333 ( .B(n4406), .A(n4405), .Z(n4407) );
  CND3X1 U2334 ( .A(n4053), .B(n4054), .C(n4063), .Z(n4024) );
  CAN2X1 U2335 ( .A(res_not_wire[48]), .B(n3841), .Z(n3447) );
  CNR2IX1 U2336 ( .B(n3422), .A(n3788), .Z(n3871) );
  CND2X1 U2337 ( .A(n3821), .B(n3450), .Z(n3788) );
  CNIVX1 U2338 ( .A(n4476), .Z(n3320) );
  CND2X1 U2339 ( .A(n3475), .B(n3765), .Z(n4503) );
  CND2X1 U2340 ( .A(n3349), .B(n3198), .Z(n3599) );
  CND2X1 U2341 ( .A(n4098), .B(n3443), .Z(n4152) );
  CENX1 U2342 ( .A(opera2[11]), .B(n3197), .Z(n4151) );
  CENX1 U2343 ( .A(opera2[12]), .B(n3197), .Z(n4188) );
  CENX1 U2344 ( .A(opera2[16]), .B(n3195), .Z(n4197) );
  CENX1 U2345 ( .A(opera2[13]), .B(n3197), .Z(n4271) );
  CENX1 U2346 ( .A(opera2[15]), .B(n3197), .Z(n4313) );
  CNR3XL U2347 ( .A(n4115), .B(n4120), .C(n4336), .Z(n4113) );
  CNR2IX1 U2348 ( .B(res_not_wire[26]), .A(n3229), .Z(n3589) );
  CNR2IX1 U2349 ( .B(n4304), .A(n4222), .Z(n3590) );
  CENX1 U2350 ( .A(opera2[19]), .B(n3195), .Z(n4371) );
  CND2X1 U2351 ( .A(n3545), .B(n3432), .Z(n3543) );
  CND2X1 U2352 ( .A(n3341), .B(n3342), .Z(n3981) );
  COND1XL U2353 ( .A(n3756), .B(n3437), .C(n3755), .Z(n3339) );
  CND2X1 U2354 ( .A(n4394), .B(n4495), .Z(n3497) );
  CND4X1 U2355 ( .A(n3227), .B(n3438), .C(i[6]), .D(i[7]), .Z(n4569) );
  CND2X1 U2356 ( .A(n3289), .B(n4079), .Z(n3611) );
  CANR2X1 U2357 ( .A(n3987), .B(n3986), .C(n3985), .D(n3984), .Z(n3993) );
  CEOX1 U2358 ( .A(result[60]), .B(n3748), .Z(n3994) );
  CND2IX1 U2359 ( .B(n4052), .A(n4024), .Z(n4041) );
  CENX1 U2360 ( .A(n3442), .B(n3728), .Z(n3441) );
  CENX1 U2361 ( .A(n4145), .B(n3312), .Z(n4146) );
  CENX1 U2362 ( .A(n3443), .B(n3327), .Z(n4183) );
  CNIVXL U2363 ( .A(n4261), .Z(n3327) );
  CNIVXL U2364 ( .A(n4314), .Z(n3312) );
  CENX1 U2365 ( .A(n1891), .B(n3377), .Z(n4279) );
  CENX1 U2366 ( .A(n3287), .B(n3197), .Z(n3318) );
  CMXI2XL U2367 ( .A0(n4625), .A1(n4623), .S(i[16]), .Z(n938) );
  CIVX3 U2368 ( .A(result[25]), .Z(n2338) );
  CNR2IX1 U2369 ( .B(n4298), .A(n4297), .Z(n4299) );
  CENX1 U2370 ( .A(res_not_wire[40]), .B(n3399), .Z(n3830) );
  CENX1 U2371 ( .A(n3925), .B(n3926), .Z(n3877) );
  COND1XL U2372 ( .A(n4076), .B(n3394), .C(n4075), .Z(n919) );
  CND3XL U2373 ( .A(n4142), .B(n4141), .C(n4140), .Z(n817) );
  CND3XL U2374 ( .A(n4361), .B(n4360), .C(n4359), .Z(n796) );
  CENX1 U2375 ( .A(n3295), .B(n3814), .Z(n3820) );
  CND2X1 U2376 ( .A(n3344), .B(n3345), .Z(n3933) );
  CMX2X1 U2377 ( .A0(n4583), .A1(n4589), .S(i[12]), .Z(n942) );
  CANR1XL U2378 ( .A(n3259), .B(n4649), .C(n4603), .Z(n4604) );
  COND1XL U2379 ( .A(n4620), .B(n4645), .C(n4619), .Z(n931) );
  COND1XL U2380 ( .A(n3306), .B(n3414), .C(n3651), .Z(n3214) );
  CAN2X1 U2381 ( .A(n3584), .B(n4392), .Z(n3217) );
  CAN3X2 U2382 ( .A(n1472), .B(n1849), .C(res_not_wire[2]), .Z(n3218) );
  COR2X1 U2383 ( .A(n3237), .B(n118), .Z(n3219) );
  CAN4X1 U2384 ( .A(i[2]), .B(i[1]), .C(i[0]), .D(i[3]), .Z(n3227) );
  CND2X1 U2385 ( .A(n3581), .B(n4512), .Z(n4385) );
  CIVX2 U2386 ( .A(n4385), .Z(n3500) );
  CAN2X1 U2387 ( .A(result[32]), .B(n4293), .Z(n3232) );
  CAN2X1 U2388 ( .A(n3455), .B(n3457), .Z(n3233) );
  CNIVXL U2389 ( .A(n4477), .Z(n3235) );
  CND2X1 U2390 ( .A(n4223), .B(n3202), .Z(n4303) );
  CND2X1 U2391 ( .A(result[0]), .B(n3500), .Z(n4553) );
  CAN2X1 U2392 ( .A(n3860), .B(n3862), .Z(n3239) );
  CND2X1 U2393 ( .A(result[53]), .B(n3649), .Z(n3849) );
  CIVXL U2394 ( .A(res_not_wire[2]), .Z(n2391) );
  CIVDXL U2395 ( .A(i[18]), .Z0(n3259), .Z1(n3260) );
  CND3XL U2396 ( .A(n4258), .B(n4257), .C(n4256), .Z(n820) );
  CNIVX1 U2397 ( .A(n820), .Z(n3261) );
  CNIVX1 U2398 ( .A(n954), .Z(n3262) );
  CNIVXL U2399 ( .A(n886), .Z(n3263) );
  CNIVX1 U2400 ( .A(n2382), .Z(n3264) );
  CNIVX1 U2401 ( .A(n952), .Z(n3265) );
  CMXI2XL U2402 ( .A0(n4600), .A1(n4601), .S(n3259), .Z(n936) );
  CNIVX1 U2403 ( .A(i[19]), .Z(n3266) );
  CNIVX1 U2404 ( .A(n928), .Z(n3267) );
  CNIVX1 U2405 ( .A(n925), .Z(n3268) );
  CNIVXL U2406 ( .A(muordi), .Z(n3291) );
  CNIVX1 U2407 ( .A(n3289), .Z(n3269) );
  CND3X1 U2408 ( .A(n4207), .B(n4206), .C(n4205), .Z(n801) );
  CENXL U2409 ( .A(opera2[24]), .B(n3197), .Z(n4203) );
  CNIVX1 U2410 ( .A(n806), .Z(n3270) );
  COND3X1 U2411 ( .A(n4379), .B(n3394), .C(n4378), .D(n4377), .Z(n806) );
  CNIVX1 U2412 ( .A(n3318), .Z(n3271) );
  CNIVX1 U2413 ( .A(n4351), .Z(n3272) );
  CENXL U2414 ( .A(opera2[29]), .B(n3197), .Z(n4351) );
  CNIVX1 U2415 ( .A(n4349), .Z(n3273) );
  COND3X1 U2416 ( .A(n4350), .B(n3212), .C(n3273), .D(n4348), .Z(n798) );
  CENXL U2417 ( .A(opera2[21]), .B(n3195), .Z(n4335) );
  CND2X1 U2418 ( .A(n4375), .B(n4328), .Z(n4331) );
  CEOXL U2419 ( .A(opera2[17]), .B(n3197), .Z(n3455) );
  CNIVX1 U2420 ( .A(n810), .Z(n3274) );
  CENXL U2421 ( .A(opera2[23]), .B(n3197), .Z(n4306) );
  CNIVX1 U2422 ( .A(n812), .Z(n3275) );
  CNIVX1 U2423 ( .A(n816), .Z(n3276) );
  CNIVX1 U2424 ( .A(n824), .Z(n3277) );
  CIVDX1 U2425 ( .A(n4352), .Z0(n4286) );
  CENXL U2426 ( .A(opera2[28]), .B(n3197), .Z(n4352) );
  COND3X2 U2427 ( .A(n4202), .B(n3212), .C(n4201), .D(n4200), .Z(n809) );
  CNIVX1 U2428 ( .A(n813), .Z(n3279) );
  CNIVX1 U2429 ( .A(n819), .Z(n3280) );
  CNIVX1 U2430 ( .A(n823), .Z(n3281) );
  CNIVX1 U2431 ( .A(n814), .Z(n3282) );
  CENXL U2432 ( .A(opera2[20]), .B(n3197), .Z(n4336) );
  CNIVX1 U2433 ( .A(n822), .Z(n3283) );
  CNIVX1 U2434 ( .A(n3285), .Z(n3284) );
  CNIVX1 U2435 ( .A(n825), .Z(n3285) );
  CIVXL U2436 ( .A(res_not_wire[0]), .Z(n2393) );
  CNIVX1 U2437 ( .A(opera2[31]), .Z(n3286) );
  CNIVX1 U2438 ( .A(opera2[30]), .Z(n3287) );
  CEOXL U2439 ( .A(n3286), .B(n3287), .Z(n4289) );
  COND2XL U2440 ( .A(n4585), .B(n3374), .C(n4586), .D(n3373), .Z(n946) );
  CMXI2X2 U2441 ( .A0(n4643), .A1(n3411), .S(i[28]), .Z(n926) );
  CMXI2X2 U2442 ( .A0(n4581), .A1(n4580), .S(i[11]), .Z(n943) );
  CDLY1XL U2443 ( .A(start), .Z(n3288) );
  CANR2XL U2444 ( .A(n3508), .B(n2347), .C(result[31]), .D(n3503), .Z(n2568)
         );
  CMXI2XL U2445 ( .A0(n3612), .A1(n3541), .S(n3611), .Z(n956) );
  CNIVX1 U2446 ( .A(n4654), .Z(n3289) );
  CNIVX1 U2447 ( .A(n956), .Z(n3290) );
  CND2IX2 U2448 ( .B(i[31]), .A(n3539), .Z(n3542) );
  CIVX1 U2449 ( .A(n4642), .Z(n3551) );
  CND2X1 U2450 ( .A(result[58]), .B(n3758), .Z(n4402) );
  CND2X1 U2451 ( .A(result[58]), .B(n3758), .Z(n3341) );
  CND2IXL U2452 ( .B(n3605), .A(n3604), .Z(n852) );
  CAN2X1 U2453 ( .A(n3403), .B(n4408), .Z(n3380) );
  CNIVX1 U2454 ( .A(n3492), .Z(n3293) );
  COND1X1 U2455 ( .A(n3430), .B(n4028), .C(n3485), .Z(n3294) );
  CIVX2 U2456 ( .A(n3468), .Z(n3295) );
  COND1X1 U2457 ( .A(n3430), .B(n4028), .C(n3485), .Z(n4404) );
  CENX1 U2458 ( .A(n3431), .B(result[56]), .Z(n3430) );
  CENX1 U2459 ( .A(n1126), .B(n4045), .Z(n3796) );
  CND2X1 U2460 ( .A(n3494), .B(n3656), .Z(n3774) );
  CND2X1 U2461 ( .A(n3473), .B(n3474), .Z(n4428) );
  CENXL U2462 ( .A(n4467), .B(n4466), .Z(n4468) );
  CND2IX1 U2463 ( .B(n3299), .A(n3643), .Z(n3965) );
  COND3XL U2464 ( .A(n4214), .B(n4384), .C(n4213), .D(n4212), .Z(n797) );
  CENX1 U2465 ( .A(result[36]), .B(n3228), .Z(n4431) );
  COND3XL U2466 ( .A(n3776), .B(n3775), .C(n3205), .D(n3831), .Z(n3301) );
  CND2X1 U2467 ( .A(n3367), .B(n3351), .Z(n3729) );
  CIVX1 U2468 ( .A(n3980), .Z(n4410) );
  CIVXL U2469 ( .A(n3682), .Z(n3701) );
  CND2X1 U2470 ( .A(n3648), .B(n3647), .Z(n3777) );
  CAN2X1 U2471 ( .A(n3660), .B(n3416), .Z(n3303) );
  COR2XL U2472 ( .A(n3439), .B(n3569), .Z(n4441) );
  CIVX2 U2473 ( .A(n3368), .Z(n3304) );
  CIVX1 U2474 ( .A(n3806), .Z(n3807) );
  CND2X1 U2475 ( .A(result[50]), .B(n3643), .Z(n3305) );
  CIVXL U2476 ( .A(n3823), .Z(n4518) );
  CND2X1 U2477 ( .A(n3859), .B(n3694), .Z(n3864) );
  CIVX2 U2478 ( .A(n3644), .Z(n3645) );
  CIVX2 U2479 ( .A(n3663), .Z(n3618) );
  CND2IX1 U2480 ( .B(n3308), .A(n3650), .Z(n3640) );
  CND2X1 U2481 ( .A(n3428), .B(n3429), .Z(n3308) );
  CND2X1 U2482 ( .A(n3753), .B(n3435), .Z(n3638) );
  CIVX2 U2483 ( .A(n3640), .Z(n3753) );
  CIVX2 U2484 ( .A(n4314), .Z(n3309) );
  CIVXL U2485 ( .A(n3673), .Z(n3310) );
  CND2X1 U2486 ( .A(n3751), .B(n3750), .Z(n3752) );
  CND2X1 U2487 ( .A(result[61]), .B(n3629), .Z(n3363) );
  CND2X2 U2488 ( .A(n3731), .B(n3943), .Z(n3799) );
  CIVX1 U2489 ( .A(n3822), .Z(n4460) );
  CND2X1 U2490 ( .A(n3767), .B(n4475), .Z(n3689) );
  COND1X2 U2491 ( .A(n4022), .B(n4021), .C(n4023), .Z(n4033) );
  CIVDXL U2492 ( .A(n4327), .Z0(n3315), .Z1(n3314) );
  CND2X1 U2493 ( .A(n3369), .B(n3316), .Z(n3783) );
  CIVX1 U2494 ( .A(n3683), .Z(n3616) );
  CND2X2 U2495 ( .A(n3754), .B(n3753), .Z(n3760) );
  CND4X1 U2496 ( .A(n3534), .B(n3533), .C(n3532), .D(n3537), .Z(n3535) );
  CIVX2 U2497 ( .A(n4003), .Z(n3979) );
  CND3X1 U2498 ( .A(n3738), .B(n3799), .C(n3800), .Z(n3739) );
  CAN2X1 U2499 ( .A(n3768), .B(n3769), .Z(n3398) );
  CIVX2 U2500 ( .A(n3836), .Z(n3776) );
  CND2X1 U2501 ( .A(n3725), .B(n3724), .Z(n3822) );
  CND2IX1 U2502 ( .B(n4398), .A(n3294), .Z(n4002) );
  CIVX2 U2503 ( .A(n3698), .Z(n3317) );
  CMXI2XL U2504 ( .A0(n4289), .A1(n4290), .S(n4362), .Z(n4301) );
  CND2X2 U2505 ( .A(n4032), .B(n4033), .Z(n4034) );
  COND3X4 U2506 ( .A(n3571), .B(n4443), .C(n4440), .D(n4442), .Z(n4447) );
  CND2X1 U2507 ( .A(n4475), .B(n3326), .Z(n4484) );
  CND2X1 U2508 ( .A(n3369), .B(n3782), .Z(n3784) );
  CIVX2 U2509 ( .A(n3755), .Z(n3624) );
  CENX1 U2510 ( .A(n3271), .B(n4362), .Z(n4369) );
  CND2IXL U2511 ( .B(n4224), .A(n4338), .Z(n4225) );
  CNR2IX1 U2512 ( .B(result[59]), .A(n3501), .Z(n4412) );
  CANR2XL U2513 ( .A(n3506), .B(n2380), .C(result[59]), .D(n3503), .Z(n2596)
         );
  CND2X1 U2514 ( .A(n3838), .B(n3338), .Z(n3319) );
  CND2XL U2515 ( .A(n3323), .B(result[42]), .Z(n3860) );
  CND3X1 U2516 ( .A(n3369), .B(n4418), .C(n3762), .Z(n3785) );
  COR2XL U2517 ( .A(n4625), .B(n4607), .Z(n4601) );
  COAN1XL U2518 ( .A(n4645), .B(i[16]), .C(n4623), .Z(n3454) );
  CND2IX1 U2519 ( .B(i[16]), .A(n4653), .Z(n3515) );
  CND2X1 U2520 ( .A(i[17]), .B(i[16]), .Z(n4607) );
  CIVX2 U2521 ( .A(n3697), .Z(n3710) );
  CND2X1 U2522 ( .A(n3618), .B(n3206), .Z(n3695) );
  CIVX2 U2523 ( .A(n3358), .Z(n3367) );
  CAN2X1 U2524 ( .A(n4545), .B(n4544), .Z(n4546) );
  CND2X2 U2525 ( .A(n4447), .B(n4441), .Z(n4432) );
  CIVX2 U2526 ( .A(n3832), .Z(n3834) );
  CND2X1 U2527 ( .A(n3638), .B(n3637), .Z(n3706) );
  CND2X1 U2528 ( .A(n3332), .B(n3333), .Z(n4511) );
  COND1X1 U2529 ( .A(n4382), .B(n4381), .C(n3165), .Z(n4121) );
  CIVXL U2530 ( .A(n3714), .Z(n3712) );
  CND3X1 U2531 ( .A(n4031), .B(n4030), .C(n4061), .Z(n4032) );
  CENX1 U2532 ( .A(opera1[5]), .B(opera1[31]), .Z(n3554) );
  CENX1 U2533 ( .A(opera1[24]), .B(opera1[31]), .Z(n3636) );
  CENX4 U2534 ( .A(opera1[13]), .B(opera1[31]), .Z(n3670) );
  CEOX4 U2535 ( .A(opera1[1]), .B(opera1[31]), .Z(n3452) );
  COAN1XL U2536 ( .A(n3427), .B(n3324), .C(n3760), .Z(n3484) );
  COND1X1 U2537 ( .A(n3324), .B(n3427), .C(n3760), .Z(n3761) );
  CND2X1 U2538 ( .A(n4419), .B(n4029), .Z(n4061) );
  CIVX1 U2539 ( .A(n3658), .Z(n3675) );
  CANR3X1 U2540 ( .A(n3483), .B(n3476), .C(n4047), .D(n4553), .Z(n4048) );
  CNR2X2 U2541 ( .A(n3638), .B(n3636), .Z(n3324) );
  CENXL U2542 ( .A(n3455), .B(n3314), .Z(n4328) );
  CNR2XL U2543 ( .A(n3688), .B(n3684), .Z(n3685) );
  CND2XL U2544 ( .A(n4345), .B(n4344), .Z(n4346) );
  CENXL U2545 ( .A(opera2[5]), .B(n3195), .Z(n4249) );
  CND2X2 U2546 ( .A(n3810), .B(n3988), .Z(n3361) );
  CNR3X1 U2547 ( .A(n3664), .B(n3670), .C(n3663), .Z(n3668) );
  COR2X1 U2548 ( .A(n3415), .B(n3495), .Z(n3642) );
  COND3X4 U2549 ( .A(n3776), .B(n3775), .C(n4547), .D(n3831), .Z(n3966) );
  COND1X2 U2550 ( .A(n3863), .B(n4466), .C(n3862), .Z(n3325) );
  COND1X1 U2551 ( .A(n4478), .B(n3235), .C(n3320), .Z(n3326) );
  CANR1X1 U2552 ( .A(n4531), .B(n4530), .C(n4529), .Z(n4532) );
  CNR2X1 U2553 ( .A(i[11]), .B(n3515), .Z(n3534) );
  CNR2X1 U2554 ( .A(i[11]), .B(i[19]), .Z(n3536) );
  CND2X1 U2555 ( .A(n4649), .B(n3329), .Z(n3330) );
  CND2X1 U2556 ( .A(n3330), .B(n3411), .Z(n4648) );
  CIVX2 U2557 ( .A(i[28]), .Z(n3329) );
  CND2X2 U2558 ( .A(n4653), .B(n4642), .Z(n4645) );
  CIVXL U2559 ( .A(n4648), .Z(n4646) );
  CIVX2 U2560 ( .A(n4505), .Z(n3331) );
  COAN1XL U2561 ( .A(n3398), .B(result[47]), .C(n3770), .Z(n3334) );
  COND1X1 U2562 ( .A(n4396), .B(n4003), .C(n4002), .Z(n4004) );
  CENXL U2563 ( .A(opera2[25]), .B(n3197), .Z(n4381) );
  CND3XL U2564 ( .A(n3483), .B(n3476), .C(n4061), .Z(n4064) );
  CIVX1 U2565 ( .A(n3490), .Z(n3337) );
  CENXL U2566 ( .A(n4007), .B(n4006), .Z(n4012) );
  CIVX2 U2567 ( .A(n3775), .Z(n3338) );
  CANR1X2 U2568 ( .A(n3297), .B(n3833), .C(n3319), .Z(n3805) );
  CND2X1 U2569 ( .A(n3376), .B(n3991), .Z(n3992) );
  CANR1X1 U2570 ( .A(n4005), .B(n3376), .C(n4004), .Z(n4006) );
  CNIVX1 U2571 ( .A(n4062), .Z(n3476) );
  CNR2IX1 U2572 ( .B(n4042), .A(n4044), .Z(n3376) );
  CND2X2 U2573 ( .A(n3355), .B(opera1[31]), .Z(n3357) );
  CND2X1 U2574 ( .A(n2335), .B(n3339), .Z(n3342) );
  CND2X1 U2575 ( .A(n4402), .B(n3981), .Z(n4397) );
  CANR1XL U2576 ( .A(n3487), .B(n3651), .C(n3337), .Z(n3766) );
  CND2X1 U2577 ( .A(n3927), .B(n3302), .Z(n3344) );
  CNR2X1 U2578 ( .A(n3346), .B(n3216), .Z(n3347) );
  CNR2X1 U2579 ( .A(n3347), .B(n3846), .Z(n4531) );
  CIVXL U2580 ( .A(n3849), .Z(n3346) );
  COND2XL U2581 ( .A(n4533), .B(n4025), .C(n4531), .D(n4027), .Z(n3812) );
  CAN2X1 U2582 ( .A(n3209), .B(n3425), .Z(n4482) );
  CNR2X2 U2583 ( .A(n4480), .B(n3219), .Z(n3841) );
  CND3X1 U2584 ( .A(n3741), .B(n3861), .C(n3239), .Z(n3742) );
  COND1X1 U2585 ( .A(n4553), .B(n3798), .C(n3797), .Z(n827) );
  CEOX4 U2586 ( .A(opera1[5]), .B(opera1[31]), .Z(n3351) );
  CENXL U2587 ( .A(n4493), .B(n4492), .Z(n4501) );
  CANR1X1 U2588 ( .A(n4491), .B(n4490), .C(n4489), .Z(n4492) );
  CND4XL U2589 ( .A(n3668), .B(n3206), .C(n3667), .D(n3665), .Z(n3676) );
  CNR2X2 U2590 ( .A(n3825), .B(n3802), .Z(n3801) );
  CND2X2 U2591 ( .A(n3356), .B(n3357), .Z(n3492) );
  CIVX2 U2592 ( .A(opera1[7]), .Z(n3355) );
  CND2X2 U2593 ( .A(n3469), .B(n3618), .Z(n3358) );
  CANR1X1 U2594 ( .A(n4649), .B(n3552), .C(n3551), .Z(n4623) );
  CND2XL U2595 ( .A(n3544), .B(n3540), .Z(n4392) );
  COAN1XL U2596 ( .A(n4644), .B(n4645), .C(n4642), .Z(n3411) );
  CENX1 U2597 ( .A(opera2[2]), .B(opera2_63), .Z(n4242) );
  CEOXL U2598 ( .A(opera2[18]), .B(n3195), .Z(n3457) );
  CND3X2 U2599 ( .A(n3362), .B(n3691), .C(n3491), .Z(n3692) );
  CIVX2 U2600 ( .A(n3361), .Z(n3362) );
  CIVX1 U2601 ( .A(n3692), .Z(n3741) );
  CND2IX1 U2602 ( .B(result[46]), .A(n3678), .Z(n3679) );
  CNR3X2 U2603 ( .A(n3556), .B(n3557), .C(n3555), .Z(n3666) );
  COR2XL U2604 ( .A(n4365), .B(n3815), .Z(n4422) );
  CANR3X1 U2605 ( .A(n3211), .B(n4010), .C(n4009), .D(n4008), .Z(n4011) );
  CIVXL U2606 ( .A(n4425), .Z(n3364) );
  CND2X1 U2607 ( .A(n108), .B(n3364), .Z(n3365) );
  COAN1X1 U2608 ( .A(n3563), .B(n3477), .C(n3562), .Z(n3366) );
  CIVX1 U2609 ( .A(n3565), .Z(n3563) );
  CIVX1 U2610 ( .A(n3358), .Z(n3368) );
  CND2IX1 U2611 ( .B(n4041), .A(n4047), .Z(n3369) );
  CIVX3 U2612 ( .A(n4645), .Z(n4649) );
  CIVX2 U2613 ( .A(n4384), .Z(n4375) );
  COND1X1 U2614 ( .A(n4478), .B(n3235), .C(n3320), .Z(n4490) );
  CND2IX1 U2615 ( .B(n4041), .A(n4047), .Z(n4018) );
  COND1XL U2616 ( .A(n3444), .B(c_inop1), .C(n3566), .Z(n4294) );
  CIVXL U2617 ( .A(n3708), .Z(n3702) );
  CIVX2 U2618 ( .A(n3426), .Z(n3383) );
  CIVX2 U2619 ( .A(n4059), .Z(n4049) );
  CND2X2 U2620 ( .A(c_inop1), .B(n3452), .Z(n3375) );
  CIVXL U2621 ( .A(n4516), .Z(n3948) );
  COND1X1 U2622 ( .A(n3702), .B(n3701), .C(n3700), .Z(n3703) );
  CIVX1 U2623 ( .A(n3968), .Z(n4481) );
  CIVX2 U2624 ( .A(n3811), .Z(n3382) );
  COND1XL U2625 ( .A(n3563), .B(n3477), .C(n3562), .Z(n3570) );
  CIVX2 U2626 ( .A(n4370), .Z(n4223) );
  CENXL U2627 ( .A(opera2[14]), .B(n3197), .Z(n4315) );
  CND2XL U2628 ( .A(c_inop1), .B(n3444), .Z(n3566) );
  CENXL U2629 ( .A(opera2[26]), .B(n3195), .Z(n4120) );
  CND4XL U2630 ( .A(res_not_wire[6]), .B(n3218), .C(n4176), .D(c_inres), .Z(
        n3377) );
  COR2X1 U2631 ( .A(n3378), .B(n4088), .Z(n3379) );
  CND2X2 U2632 ( .A(n3624), .B(n3623), .Z(n3751) );
  CNR2X2 U2633 ( .A(n3380), .B(n4407), .Z(n4409) );
  CIVX2 U2634 ( .A(n4409), .Z(n3426) );
  CIVX1 U2635 ( .A(n3864), .Z(n3899) );
  CNIVX1 U2636 ( .A(n4652), .Z(n3508) );
  CEOXL U2637 ( .A(n4460), .B(n4459), .Z(n3826) );
  CND2X1 U2638 ( .A(n3733), .B(n3732), .Z(n3737) );
  CND2IX1 U2639 ( .B(n3598), .A(n4439), .Z(n4430) );
  CND2X2 U2640 ( .A(n4119), .B(n4307), .Z(n4382) );
  CENX1 U2641 ( .A(result[40]), .B(n3716), .Z(n3717) );
  CANR2X1 U2642 ( .A(n3508), .B(n4656), .C(result[0]), .D(n3505), .Z(n2531) );
  CND2XL U2643 ( .A(n3886), .B(n3885), .Z(n3892) );
  CND3XL U2644 ( .A(n3211), .B(n4036), .C(n4074), .Z(n4037) );
  COND3X1 U2645 ( .A(n4527), .B(n3496), .C(n4526), .D(n4525), .Z(n849) );
  COND3X1 U2646 ( .A(n3913), .B(n3212), .C(n3912), .D(n3911), .Z(n851) );
  COND1XL U2647 ( .A(n4046), .B(res_not_wire[60]), .C(n3207), .Z(n3392) );
  CANR2XL U2648 ( .A(n3507), .B(n2361), .C(result[6]), .D(n3504), .Z(n2543) );
  CANR2XL U2649 ( .A(n3508), .B(n2338), .C(result[25]), .D(n3503), .Z(n2562)
         );
  CANR2XL U2650 ( .A(n3507), .B(n2357), .C(result[24]), .D(n3504), .Z(n2561)
         );
  CANR2XL U2651 ( .A(n3506), .B(n2367), .C(result[26]), .D(n3503), .Z(n2563)
         );
  CNR2X1 U2652 ( .A(n3968), .B(n4480), .Z(n3400) );
  CND2XL U2653 ( .A(result[32]), .B(n4293), .Z(n3914) );
  COAN1X1 U2654 ( .A(n3297), .B(n3692), .C(n3382), .Z(n3743) );
  CND2X1 U2655 ( .A(n3426), .B(n3980), .Z(n3385) );
  CIVX1 U2656 ( .A(n3401), .Z(n3501) );
  CND2XL U2657 ( .A(n4649), .B(n4631), .Z(n4625) );
  CNR2IX1 U2658 ( .B(n3207), .A(n3404), .Z(n4124) );
  CIVX1 U2659 ( .A(n4530), .Z(n3813) );
  CND2XL U2660 ( .A(n4649), .B(n4609), .Z(n4610) );
  CIVX1 U2661 ( .A(n4572), .Z(n4585) );
  CND3X1 U2662 ( .A(n3785), .B(n3784), .C(n3783), .Z(n3787) );
  COR2XL U2663 ( .A(n4448), .B(n4447), .Z(n4449) );
  CND2X1 U2664 ( .A(n3767), .B(n4479), .Z(n4488) );
  CND2X1 U2665 ( .A(n3725), .B(n3824), .Z(n3803) );
  CND2XL U2666 ( .A(n4649), .B(n4624), .Z(n4622) );
  CEOXL U2667 ( .A(n3340), .B(n3386), .Z(n4461) );
  CANR1XL U2668 ( .A(n4460), .B(n4459), .C(n4458), .Z(n3386) );
  COR2XL U2669 ( .A(n4607), .B(n4606), .Z(n4609) );
  CND2XL U2670 ( .A(n4585), .B(n4584), .Z(n4589) );
  CND2IXL U2671 ( .B(n3599), .A(n4481), .Z(n3600) );
  CNR2X2 U2672 ( .A(n3522), .B(n3521), .Z(n3530) );
  COAN1XL U2673 ( .A(n3227), .B(n4645), .C(n4642), .Z(n3407) );
  CAN3XL U2674 ( .A(n4481), .B(n3450), .C(n3412), .Z(n3409) );
  CND2IXL U2675 ( .B(n3970), .A(n3969), .Z(n3971) );
  CND2IXL U2676 ( .B(n3869), .A(n3868), .Z(n3870) );
  CIVXL U2677 ( .A(n4115), .Z(n4224) );
  CIVXL U2678 ( .A(n4440), .Z(n4446) );
  CENX2 U2679 ( .A(result[43]), .B(n3704), .Z(n4466) );
  COND1X2 U2680 ( .A(n3568), .B(n3232), .C(n3567), .Z(n3887) );
  CNR2IXL U2681 ( .B(result[39]), .A(n3501), .Z(n3950) );
  CIVXL U2682 ( .A(n4637), .Z(n4634) );
  CNR2IXL U2683 ( .B(result[56]), .A(n3501), .Z(n3816) );
  CANR2XL U2684 ( .A(n3507), .B(n2368), .C(result[20]), .D(n3504), .Z(n2557)
         );
  CANR2XL U2685 ( .A(n3507), .B(n2363), .C(result[2]), .D(n3504), .Z(n2539) );
  CANR2XL U2686 ( .A(n3507), .B(n2362), .C(result[4]), .D(n3504), .Z(n2541) );
  CANR2XL U2687 ( .A(n4652), .B(n3242), .C(result[33]), .D(n3413), .Z(n2570)
         );
  CANR2XL U2688 ( .A(n3507), .B(n2353), .C(result[1]), .D(n3504), .Z(n2538) );
  CANR2XL U2689 ( .A(n3507), .B(n2351), .C(result[5]), .D(n3504), .Z(n2542) );
  CNR2XL U2690 ( .A(n4640), .B(n2284), .Z(n4636) );
  CND2IXL U2691 ( .B(n3387), .A(n3893), .Z(n879) );
  CNR2X1 U2692 ( .A(n3255), .B(n3509), .Z(n3387) );
  CND2IXL U2693 ( .B(n3388), .A(n3937), .Z(n869) );
  CNR2X1 U2694 ( .A(n3256), .B(n3509), .Z(n3388) );
  CND2IXL U2695 ( .B(n3389), .A(n4073), .Z(n867) );
  CNR2X1 U2696 ( .A(n3257), .B(n3509), .Z(n3389) );
  CND2IXL U2697 ( .B(n3390), .A(n4555), .Z(n864) );
  CNR2X1 U2698 ( .A(n3252), .B(n3509), .Z(n3390) );
  CND2IX1 U2699 ( .B(n3391), .A(n3936), .Z(n881) );
  CNR2X1 U2700 ( .A(n3258), .B(n3509), .Z(n3391) );
  CND2XL U2701 ( .A(n3502), .B(n3914), .Z(n3917) );
  CND2XL U2702 ( .A(n3502), .B(n4433), .Z(n4436) );
  CANR2XL U2703 ( .A(n3506), .B(n2327), .C(result[51]), .D(n3503), .Z(n2588)
         );
  CNR2IXL U2704 ( .B(result[48]), .A(n3501), .Z(n4496) );
  CANR2XL U2705 ( .A(n3508), .B(n3442), .C(result[37]), .D(n3503), .Z(n2574)
         );
  CANR2XL U2706 ( .A(n3507), .B(n2343), .C(result[21]), .D(n3504), .Z(n2558)
         );
  CANR2XL U2707 ( .A(n3507), .B(n2339), .C(result[19]), .D(n3504), .Z(n2556)
         );
  CANR2XL U2708 ( .A(n3506), .B(n3321), .C(result[48]), .D(n3503), .Z(n2585)
         );
  CANR2XL U2709 ( .A(n3508), .B(n3249), .C(result[39]), .D(n3503), .Z(n2576)
         );
  CANR2XL U2710 ( .A(n3507), .B(n2346), .C(result[23]), .D(n3504), .Z(n2560)
         );
  CANR2XL U2711 ( .A(n3506), .B(n3221), .C(result[44]), .D(n3503), .Z(n2581)
         );
  CANR2XL U2712 ( .A(n3506), .B(n2354), .C(result[22]), .D(n3504), .Z(n2559)
         );
  CNR2IXL U2713 ( .B(result[55]), .A(n3501), .Z(n4535) );
  CND2IXL U2714 ( .B(n4384), .A(n4308), .Z(n4311) );
  CND2XL U2715 ( .A(n3502), .B(n3888), .Z(n3891) );
  CND2XL U2716 ( .A(n4375), .B(n4146), .Z(n4149) );
  CND2XL U2717 ( .A(n4375), .B(n4162), .Z(n4165) );
  CND2XL U2718 ( .A(n4375), .B(n3166), .Z(n4172) );
  CND2XL U2719 ( .A(n4375), .B(n4183), .Z(n4186) );
  CND2XL U2720 ( .A(n4375), .B(n4281), .Z(n4284) );
  CEOX1 U2721 ( .A(n1476), .B(n4074), .Z(n4076) );
  CND2IXL U2722 ( .B(n4660), .A(n3200), .Z(n4075) );
  CNR2IXL U2723 ( .B(result[57]), .A(n3501), .Z(n4423) );
  CNR2IXL U2724 ( .B(result[29]), .A(n3499), .Z(n4211) );
  CNR2IXL U2725 ( .B(result[23]), .A(n3498), .Z(n4227) );
  CNR2IXL U2726 ( .B(result[54]), .A(n3501), .Z(n3855) );
  CNR2IXL U2727 ( .B(result[36]), .A(n3501), .Z(n4434) );
  CNR2IXL U2728 ( .B(result[35]), .A(n3501), .Z(n4451) );
  CNR2IXL U2729 ( .B(result[40]), .A(n3501), .Z(n4524) );
  CNR2IXL U2730 ( .B(result[50]), .A(n3501), .Z(n4550) );
  CNR2IXL U2731 ( .B(result[52]), .A(n3501), .Z(n4508) );
  CNR2IXL U2732 ( .B(result[41]), .A(n3501), .Z(n3827) );
  CNR2IXL U2733 ( .B(result[45]), .A(n3501), .Z(n3874) );
  CNR2IXL U2734 ( .B(result[53]), .A(n3501), .Z(n3881) );
  CNR2IXL U2735 ( .B(result[38]), .A(n3501), .Z(n3910) );
  CNR2IXL U2736 ( .B(result[51]), .A(n3501), .Z(n3975) );
  CNR2IXL U2737 ( .B(result[63]), .A(n3501), .Z(n4035) );
  CNR2IXL U2738 ( .B(result[42]), .A(n3501), .Z(n4462) );
  CNR2IXL U2739 ( .B(result[43]), .A(n3501), .Z(n4470) );
  CNR2IXL U2740 ( .B(result[49]), .A(n3501), .Z(n3842) );
  CNR2IXL U2741 ( .B(result[34]), .A(n3501), .Z(n3889) );
  CNR2IXL U2742 ( .B(result[22]), .A(n3498), .Z(n4339) );
  CNR2IXL U2743 ( .B(result[28]), .A(n3498), .Z(n4347) );
  CNR2IXL U2744 ( .B(result[7]), .A(n3498), .Z(n4178) );
  CNR2IXL U2745 ( .B(result[11]), .A(n3499), .Z(n4184) );
  CNR2IXL U2746 ( .B(result[13]), .A(n3498), .Z(n4193) );
  CNR2IXL U2747 ( .B(result[2]), .A(n3498), .Z(n4236) );
  CNR2IXL U2748 ( .B(result[6]), .A(n3499), .Z(n4255) );
  CNR2IXL U2749 ( .B(result[10]), .A(n3498), .Z(n4265) );
  CNR2IXL U2750 ( .B(result[14]), .A(n3498), .Z(n4274) );
  CNR2IXL U2751 ( .B(result[8]), .A(n3498), .Z(n4282) );
  CNR2IXL U2752 ( .B(result[24]), .A(n3498), .Z(n4309) );
  CNR2IXL U2753 ( .B(result[16]), .A(n3498), .Z(n4320) );
  CNR2IXL U2754 ( .B(result[18]), .A(n3498), .Z(n4329) );
  COAN1XL U2755 ( .A(n4645), .B(i[0]), .C(n4642), .Z(n3453) );
  CANR2XL U2756 ( .A(n3507), .B(n2352), .C(result[3]), .D(n3504), .Z(n2540) );
  CNR2IX1 U2757 ( .B(i[2]), .A(n4562), .Z(n3959) );
  CMX2XL U2758 ( .A0(n3420), .A1(n4618), .S(i[22]), .Z(n932) );
  CMX2XL U2759 ( .A0(n3418), .A1(n4566), .S(i[6]), .Z(n948) );
  CMX2XL U2760 ( .A0(n4621), .A1(n4627), .S(i[24]), .Z(n930) );
  CNR2IXL U2761 ( .B(result[19]), .A(n3498), .Z(n4219) );
  CMXI2XL U2762 ( .A0(n3508), .A1(n3505), .S(result[35]), .Z(n3894) );
  CMXI2XL U2763 ( .A0(n3508), .A1(n3505), .S(result[36]), .Z(n3906) );
  CMXI2XL U2764 ( .A0(n3508), .A1(n3505), .S(result[49]), .Z(n3955) );
  CMXI2XL U2765 ( .A0(n3508), .A1(n3505), .S(result[43]), .Z(n4071) );
  CNR2IXL U2766 ( .B(n3234), .A(n3510), .Z(n4078) );
  CMXI2XL U2767 ( .A0(n3508), .A1(n3505), .S(result[41]), .Z(n4077) );
  CNR2IXL U2768 ( .B(res_not_wire[6]), .A(n3510), .Z(n3606) );
  CNR2IXL U2769 ( .B(n38), .A(n3510), .Z(n4557) );
  CNR2IXL U2770 ( .B(res_not_wire[24]), .A(n3510), .Z(n4558) );
  CNR2IXL U2771 ( .B(res_not_wire[26]), .A(n3510), .Z(n3613) );
  CNR2IXL U2772 ( .B(res_not_wire[42]), .A(n3510), .Z(n3897) );
  CMXI2XL U2773 ( .A0(n3508), .A1(n3505), .S(result[42]), .Z(n3896) );
  CMXI2XL U2774 ( .A0(n3508), .A1(n3505), .S(n3167), .Z(n3938) );
  CMXI2XL U2775 ( .A0(n3508), .A1(n3505), .S(result[45]), .Z(n4542) );
  CEOXL U2776 ( .A(n3286), .B(n3195), .Z(n4290) );
  CIVXL U2777 ( .A(result[56]), .Z(n2334) );
  CIVXL U2778 ( .A(result[54]), .Z(n4538) );
  CIVXL U2779 ( .A(result[47]), .Z(n4474) );
  CND2XL U2780 ( .A(n4394), .B(n4495), .Z(n3394) );
  CND2XL U2781 ( .A(n4394), .B(n4495), .Z(n3395) );
  CNR2IXL U2782 ( .B(result[46]), .A(n3501), .Z(n3930) );
  CANR2XL U2783 ( .A(n3508), .B(n2329), .C(result[46]), .D(n3503), .Z(n2583)
         );
  CIVXL U2784 ( .A(result[46]), .Z(n2329) );
  CANR1X1 U2785 ( .A(n4399), .B(n4062), .C(n4398), .Z(n4401) );
  CEOX1 U2786 ( .A(opera1[19]), .B(opera1[31]), .Z(n3397) );
  CIVXL U2787 ( .A(n3500), .Z(n3498) );
  CIVX2 U2788 ( .A(n4226), .Z(n4307) );
  CNIVX1 U2789 ( .A(n4652), .Z(n3506) );
  CND2X1 U2790 ( .A(n4649), .B(n4571), .Z(n4586) );
  CND2X1 U2791 ( .A(n4079), .B(n4495), .Z(n4384) );
  CANR1XL U2792 ( .A(n3502), .B(n4041), .C(n4040), .Z(n4070) );
  CNIVX1 U2793 ( .A(n4652), .Z(n3507) );
  CNR2IXL U2794 ( .B(n3211), .A(n4439), .Z(n3886) );
  CIVX2 U2795 ( .A(n3646), .Z(n3650) );
  CND3X1 U2796 ( .A(n3368), .B(n3303), .C(n3633), .Z(n3646) );
  CNR2IXL U2797 ( .B(n3211), .A(n3408), .Z(n4499) );
  CND2XL U2798 ( .A(n3328), .B(n3406), .Z(n4251) );
  CND2XL U2799 ( .A(n3710), .B(n3367), .Z(n3714) );
  CNR2X1 U2800 ( .A(n4537), .B(n3212), .Z(n3854) );
  CAN2XL U2801 ( .A(n4419), .B(n3781), .Z(n3782) );
  COND1XL U2802 ( .A(n3468), .B(n4403), .C(n4026), .Z(n4030) );
  CNR2X1 U2803 ( .A(n4534), .B(n3210), .Z(n4536) );
  CNR2IXL U2804 ( .B(n3211), .A(n3928), .Z(n3873) );
  CNR2IXL U2805 ( .B(n3211), .A(n4506), .Z(n3974) );
  CNR2IXL U2806 ( .B(n3211), .A(n3409), .Z(n4456) );
  CNR2IXL U2807 ( .B(n3211), .A(n3402), .Z(n3603) );
  CNR2IXL U2808 ( .B(n3502), .A(n4478), .Z(n3903) );
  CAN2XL U2809 ( .A(n4481), .B(n3412), .Z(n3399) );
  CAN2X1 U2810 ( .A(n4656), .B(n3500), .Z(n3401) );
  CNR3X1 U2811 ( .A(n3217), .B(n3541), .C(n3543), .Z(n4652) );
  COND1XL U2812 ( .A(n3834), .B(n3833), .C(n3297), .Z(n3837) );
  CND2XL U2813 ( .A(n4394), .B(n4495), .Z(n3496) );
  CND2IX1 U2814 ( .B(n3630), .A(n3488), .Z(n3632) );
  CENX1 U2815 ( .A(n4307), .B(n4306), .Z(n4308) );
  CND2IX1 U2816 ( .B(n4222), .A(n4223), .Z(n4302) );
  CNR2IXL U2817 ( .B(n4519), .A(n4518), .Z(n4521) );
  COND1XL U2818 ( .A(n4518), .B(n3825), .C(n3824), .Z(n4459) );
  CNR2IX1 U2819 ( .B(n3920), .A(n3919), .Z(n3921) );
  CENX1 U2820 ( .A(n3423), .B(n3908), .Z(n3909) );
  CNIVX1 U2821 ( .A(n3413), .Z(n3505) );
  COND1XL U2822 ( .A(n4306), .B(n4226), .C(n4203), .Z(n4204) );
  CNR2X1 U2823 ( .A(n4306), .B(n4381), .Z(n4114) );
  CNR2X1 U2824 ( .A(n4335), .B(n4203), .Z(n4112) );
  CNR2X1 U2825 ( .A(n4056), .B(n4055), .Z(n4060) );
  CND2XL U2826 ( .A(n4053), .B(n4052), .Z(n4056) );
  CNR3X2 U2827 ( .A(n4242), .B(n4241), .C(n4134), .Z(n4095) );
  CANR11XL U2828 ( .A(n3209), .B(n4425), .C(n4424), .D(n4423), .Z(n4427) );
  CNR2X1 U2829 ( .A(n3593), .B(n3378), .Z(n3596) );
  CNR2X1 U2830 ( .A(n4088), .B(n3594), .Z(n3595) );
  CAN2XL U2831 ( .A(n3821), .B(n4481), .Z(n3402) );
  CND3X1 U2832 ( .A(n3310), .B(n3675), .C(n3674), .Z(n3687) );
  CND2XL U2833 ( .A(n4134), .B(n4135), .Z(n4136) );
  CND3XL U2834 ( .A(n4053), .B(n3502), .C(n3201), .Z(n4043) );
  COR2X1 U2835 ( .A(n4191), .B(n3379), .Z(n4318) );
  CANR3XL U2836 ( .A(n3999), .B(n3998), .C(n3997), .D(n3996), .Z(n4000) );
  COND1XL U2837 ( .A(n4411), .B(n3250), .C(n3222), .Z(n3998) );
  CNIVX1 U2838 ( .A(n3413), .Z(n3504) );
  CNR2X1 U2839 ( .A(n4306), .B(n4203), .Z(n4119) );
  CND2XL U2840 ( .A(n4642), .B(n4570), .Z(n4572) );
  CND2XL U2841 ( .A(n4649), .B(n4569), .Z(n4570) );
  CND2X1 U2842 ( .A(n4585), .B(n4576), .Z(n4579) );
  CND2XL U2843 ( .A(n4649), .B(n4575), .Z(n4576) );
  CND2X1 U2844 ( .A(n3415), .B(n3414), .Z(n3630) );
  CANR1X2 U2845 ( .A(n3737), .B(n3736), .C(n3735), .Z(n3800) );
  CND2XL U2846 ( .A(n4649), .B(n4588), .Z(n4584) );
  CND2XL U2847 ( .A(n4042), .B(n3988), .Z(n4027) );
  CNR2IXL U2848 ( .B(n3220), .A(n3968), .Z(n3868) );
  CNR2IXL U2849 ( .B(n3226), .A(n3968), .Z(n3969) );
  CNIVX1 U2850 ( .A(n3413), .Z(n3503) );
  CND2XL U2851 ( .A(n3727), .B(n3733), .Z(n3944) );
  CND2X1 U2852 ( .A(n4020), .B(n4019), .Z(n4023) );
  CAN2XL U2853 ( .A(n3436), .B(n4642), .Z(n3405) );
  COR2X1 U2854 ( .A(n4575), .B(n4586), .Z(n4578) );
  CND2XL U2855 ( .A(n3947), .B(n3946), .Z(n4516) );
  COND1XL U2856 ( .A(n3945), .B(n3944), .C(n3943), .Z(n3946) );
  CND2XL U2857 ( .A(n3831), .B(n4545), .Z(n3839) );
  CND2XL U2858 ( .A(n4392), .B(n4395), .Z(n921) );
  CND2X1 U2859 ( .A(n3676), .B(n3671), .Z(n3681) );
  CND2XL U2860 ( .A(n4058), .B(n4057), .Z(n4040) );
  CNR2XL U2861 ( .A(n4241), .B(n4280), .Z(n4133) );
  COND1XL U2862 ( .A(n4231), .B(n3203), .C(n2391), .Z(n4160) );
  CND2XL U2863 ( .A(n3438), .B(n3227), .Z(n4564) );
  CND2XL U2864 ( .A(n4443), .B(n4442), .Z(n4445) );
  COND1XL U2865 ( .A(n4243), .B(n4242), .C(n4241), .Z(n4244) );
  CENX1 U2866 ( .A(n1475), .B(n4269), .Z(n4270) );
  CND2XL U2867 ( .A(n4649), .B(n4633), .Z(n4635) );
  CENX1 U2868 ( .A(opera1[17]), .B(opera1[31]), .Z(n3654) );
  CANR2X1 U2869 ( .A(n4017), .B(n3354), .C(result[62]), .D(n4016), .Z(n4019)
         );
  CND2X1 U2870 ( .A(n4014), .B(n4013), .Z(n4017) );
  CANR1XL U2871 ( .A(result[45]), .B(n3200), .C(n3930), .Z(n3931) );
  CND2X1 U2872 ( .A(n3526), .B(n3525), .Z(n3527) );
  CND2XL U2873 ( .A(i[7]), .B(n4566), .Z(n4567) );
  CNR2XL U2874 ( .A(n4564), .B(i[7]), .Z(n4565) );
  CND2XL U2875 ( .A(i[15]), .B(n4596), .Z(n4597) );
  CNR2XL U2876 ( .A(n4594), .B(i[15]), .Z(n4595) );
  CND2XL U2877 ( .A(i[23]), .B(n4618), .Z(n4619) );
  CNR2XL U2878 ( .A(n4616), .B(i[23]), .Z(n4617) );
  CND2XL U2879 ( .A(i[27]), .B(n4637), .Z(n4638) );
  CNR2X1 U2880 ( .A(n4641), .B(n4640), .Z(n4644) );
  COND1X1 U2881 ( .A(n3398), .B(result[47]), .C(n3770), .Z(n4479) );
  CND3XL U2882 ( .A(result[47]), .B(n3769), .C(n3768), .Z(n3770) );
  COND2XL U2883 ( .A(i[29]), .B(n4647), .C(n4646), .D(n2281), .Z(n925) );
  CEOX1 U2884 ( .A(opera1[19]), .B(opera1[31]), .Z(n3414) );
  CEOX1 U2885 ( .A(opera1[16]), .B(n3215), .Z(n3416) );
  CEOX1 U2886 ( .A(opera2[9]), .B(opera2_63), .Z(n3417) );
  CAN2XL U2887 ( .A(n4649), .B(n4563), .Z(n3418) );
  CAN2XL U2888 ( .A(n4649), .B(n4593), .Z(n3419) );
  CAN2XL U2889 ( .A(n4649), .B(n4615), .Z(n3420) );
  CND2X1 U2890 ( .A(n3260), .B(n4602), .Z(n4605) );
  CANR1XL U2891 ( .A(n2281), .B(n4649), .C(n4648), .Z(n4650) );
  CND2XL U2892 ( .A(n4649), .B(n3227), .Z(n3957) );
  CND2XL U2893 ( .A(i[0]), .B(n4649), .Z(n4561) );
  CANR1XL U2894 ( .A(n3374), .B(n4649), .C(n4572), .Z(n4573) );
  CANR1XL U2895 ( .A(n2298), .B(n4649), .C(n4579), .Z(n4580) );
  CNR2IX1 U2896 ( .B(n4590), .A(n4589), .Z(n4591) );
  CNR2IXL U2897 ( .B(i[12]), .A(n4586), .Z(n4587) );
  CNR2IX1 U2898 ( .B(n4612), .A(n4611), .Z(n4613) );
  CNR2IX1 U2899 ( .B(n4628), .A(n4627), .Z(n4629) );
  CND2XL U2900 ( .A(n4649), .B(n4644), .Z(n4643) );
  CND2X1 U2901 ( .A(n4632), .B(n3579), .Z(n3580) );
  CNR3XL U2902 ( .A(n3578), .B(n3577), .C(n3576), .Z(n3579) );
  CND3XL U2903 ( .A(i[29]), .B(i[30]), .C(i[24]), .Z(n3577) );
  CANR1XL U2904 ( .A(result[40]), .B(n3200), .C(n3827), .Z(n3828) );
  CANR1XL U2905 ( .A(result[35]), .B(n3200), .C(n4434), .Z(n4435) );
  CND3XL U2906 ( .A(n3502), .B(n4450), .C(n4449), .Z(n4453) );
  CANR1XL U2907 ( .A(result[34]), .B(n3200), .C(n4451), .Z(n4452) );
  CENX1 U2908 ( .A(n3396), .B(n4439), .Z(n4454) );
  CANR1XL U2909 ( .A(n3940), .B(n3402), .C(res_not_wire[38]), .Z(n3954) );
  CENX1 U2910 ( .A(n4324), .B(n3241), .Z(n4202) );
  CANR1XL U2911 ( .A(result[16]), .B(n3200), .C(n4199), .Z(n4200) );
  CANR1XL U2912 ( .A(result[53]), .B(n3200), .C(n3855), .Z(n3856) );
  CANR1XL U2913 ( .A(result[62]), .B(n3200), .C(n4035), .Z(n4038) );
  CANR1XL U2914 ( .A(result[25]), .B(n3200), .C(n4386), .Z(n4387) );
  CANR1XL U2915 ( .A(result[30]), .B(n3200), .C(n4366), .Z(n4367) );
  CANR1XL U2916 ( .A(result[28]), .B(n3200), .C(n4211), .Z(n4212) );
  CANR1XL U2917 ( .A(result[22]), .B(n3200), .C(n4227), .Z(n4228) );
  CND3XL U2918 ( .A(n4375), .B(n4226), .C(n4225), .Z(n4229) );
  CNR2IX2 U2919 ( .B(n3421), .A(n4411), .Z(n4046) );
  COND1XL U2920 ( .A(n4370), .B(n146), .C(n4091), .Z(n4092) );
  COND1XL U2921 ( .A(n3968), .B(n3350), .C(n132), .Z(n3885) );
  CANR1XL U2922 ( .A(result[38]), .B(n3200), .C(n3950), .Z(n3951) );
  CNR2X1 U2923 ( .A(n3851), .B(n4658), .Z(n3791) );
  CNR2X1 U2924 ( .A(n3790), .B(n3853), .Z(n3792) );
  CND2X1 U2925 ( .A(res_not_wire[50]), .B(n3226), .Z(n3790) );
  COND1XL U2926 ( .A(n4045), .B(n3251), .C(n3223), .Z(n4036) );
  COND1XL U2927 ( .A(n4422), .B(n3252), .C(n3224), .Z(n4424) );
  CEOX1 U2928 ( .A(n3879), .B(res_not_wire[52]), .Z(n3880) );
  CEOXL U2929 ( .A(n4357), .B(res_not_wire[28]), .Z(n4210) );
  CANR1XL U2930 ( .A(result[23]), .B(n3200), .C(n4309), .Z(n4310) );
  CND2IX1 U2931 ( .B(result[49]), .A(n3774), .Z(n3831) );
  CANR1XL U2932 ( .A(result[51]), .B(n3200), .C(n4508), .Z(n4509) );
  CANR1XL U2933 ( .A(result[37]), .B(n3200), .C(n3910), .Z(n3911) );
  CANR1XL U2934 ( .A(result[39]), .B(n3200), .C(n4524), .Z(n4525) );
  COND3X1 U2935 ( .A(n4554), .B(n4553), .C(n4552), .D(n4551), .Z(n839) );
  CANR1XL U2936 ( .A(result[49]), .B(n3200), .C(n4550), .Z(n4551) );
  COND3X1 U2937 ( .A(n3884), .B(n4553), .C(n3883), .D(n3882), .Z(n836) );
  CANR1XL U2938 ( .A(result[52]), .B(n3200), .C(n3881), .Z(n3882) );
  COND3X1 U2939 ( .A(n3978), .B(n4553), .C(n3977), .D(n3976), .Z(n838) );
  CANR1XL U2940 ( .A(result[50]), .B(n3200), .C(n3975), .Z(n3976) );
  COND3X1 U2941 ( .A(n3877), .B(n4553), .C(n3876), .D(n3875), .Z(n844) );
  CANR1XL U2942 ( .A(result[44]), .B(n3200), .C(n3874), .Z(n3875) );
  CANR1XL U2943 ( .A(result[19]), .B(n3200), .C(n4376), .Z(n4377) );
  CANR1XL U2944 ( .A(result[27]), .B(n3200), .C(n4347), .Z(n4348) );
  COND3X1 U2945 ( .A(n4342), .B(n3210), .C(n4341), .D(n4340), .Z(n804) );
  CND3XL U2946 ( .A(n4375), .B(n4338), .C(n4337), .Z(n4341) );
  CANR1XL U2947 ( .A(result[21]), .B(n3200), .C(n4339), .Z(n4340) );
  CND3XL U2948 ( .A(i[28]), .B(n4649), .C(n4644), .Z(n4647) );
  CANR3X1 U2949 ( .A(n4499), .B(n4498), .C(n4497), .D(n4496), .Z(n4500) );
  CENX1 U2950 ( .A(n3787), .B(n4020), .Z(n3798) );
  CNR2IX1 U2951 ( .B(result[62]), .A(n3501), .Z(n3794) );
  CNR2IX1 U2952 ( .B(result[60]), .A(n3501), .Z(n3996) );
  CNR2IX1 U2953 ( .B(result[17]), .A(n3498), .Z(n4199) );
  CNR2IXL U2954 ( .B(result[1]), .A(n3499), .Z(n4084) );
  CNR2IXL U2955 ( .B(result[21]), .A(n3499), .Z(n4108) );
  CNR2IXL U2956 ( .B(result[27]), .A(n3498), .Z(n4126) );
  CNR2IXL U2957 ( .B(result[9]), .A(n3499), .Z(n4139) );
  CNR2IXL U2958 ( .B(result[15]), .A(n3499), .Z(n4147) );
  CNR2IXL U2959 ( .B(result[12]), .A(n3498), .Z(n4156) );
  CNR2IXL U2960 ( .B(result[3]), .A(n3499), .Z(n4163) );
  CNR2IXL U2961 ( .B(result[5]), .A(n3498), .Z(n4170) );
  CNR2IX1 U2962 ( .B(result[30]), .A(n3499), .Z(n4358) );
  CNR2IX1 U2963 ( .B(result[31]), .A(n3499), .Z(n4366) );
  CNR2IX1 U2964 ( .B(result[20]), .A(n3499), .Z(n4376) );
  CNR2IX1 U2965 ( .B(result[26]), .A(n3499), .Z(n4386) );
  CND2X1 U2966 ( .A(n3575), .B(n3574), .Z(n4624) );
  CNR2X1 U2967 ( .A(n3573), .B(n4607), .Z(n3574) );
  CNR2IXL U2968 ( .B(result[59]), .A(n4495), .Z(n3997) );
  CNR2IXL U2969 ( .B(n4661), .A(n3549), .Z(n3547) );
  CND3XL U2970 ( .A(i[1]), .B(i[0]), .C(n4649), .Z(n4562) );
  COND1XL U2971 ( .A(n3509), .B(n2408), .C(n2541), .Z(n915) );
  COND1XL U2972 ( .A(n3509), .B(n2435), .C(n2557), .Z(n899) );
  COND1XL U2973 ( .A(n128), .B(n3509), .C(n2574), .Z(n882) );
  COND1XL U2974 ( .A(n144), .B(n3510), .C(n2558), .Z(n898) );
  COND1XL U2975 ( .A(n134), .B(n3509), .C(n2568), .Z(n888) );
  COND1XL U2976 ( .A(n3509), .B(n2424), .C(n2567), .Z(n889) );
  CANR2X1 U2977 ( .A(n3508), .B(n2340), .C(result[30]), .D(n3503), .Z(n2567)
         );
  COND1XL U2978 ( .A(n146), .B(n3509), .C(n2556), .Z(n900) );
  COND1XL U2979 ( .A(n138), .B(n3509), .C(n2564), .Z(n892) );
  COND1XL U2980 ( .A(n3509), .B(n4658), .C(n2585), .Z(n871) );
  COND1XL U2981 ( .A(n3509), .B(n3237), .C(n2583), .Z(n873) );
  COND1XL U2982 ( .A(n114), .B(n3510), .C(n2588), .Z(n868) );
  COND1XL U2983 ( .A(n136), .B(n3509), .C(n2566), .Z(n890) );
  CANR2X1 U2984 ( .A(n3507), .B(n2341), .C(result[29]), .D(n3413), .Z(n2566)
         );
  COND1XL U2985 ( .A(n108), .B(n3509), .C(n2594), .Z(n862) );
  CANR2X1 U2986 ( .A(n3506), .B(n2379), .C(result[57]), .D(n3503), .Z(n2594)
         );
  COND1XL U2987 ( .A(n3510), .B(n2397), .C(n2551), .Z(n905) );
  CANR2X1 U2988 ( .A(n3507), .B(n2365), .C(result[14]), .D(n3505), .Z(n2551)
         );
  COND1XL U2989 ( .A(n3509), .B(n2396), .C(n2547), .Z(n909) );
  CANR2X1 U2990 ( .A(n3507), .B(n2360), .C(result[10]), .D(n3504), .Z(n2547)
         );
  COND1XL U2991 ( .A(n126), .B(n3509), .C(n2576), .Z(n880) );
  COND1XL U2992 ( .A(n3509), .B(n2391), .C(n2539), .Z(n917) );
  COND1XL U2993 ( .A(n142), .B(n3510), .C(n2560), .Z(n896) );
  COND1XL U2994 ( .A(n148), .B(n3510), .C(n2554), .Z(n902) );
  COND1XL U2995 ( .A(n132), .B(n3509), .C(n2570), .Z(n886) );
  COND1XL U2996 ( .A(n3509), .B(n2372), .C(n2599), .Z(n857) );
  CANR2X1 U2997 ( .A(n3506), .B(n4014), .C(result[62]), .D(n3503), .Z(n2599)
         );
  COND1XL U2998 ( .A(n3510), .B(n4657), .C(n2597), .Z(n859) );
  COND1XL U2999 ( .A(n3509), .B(n2323), .C(n2596), .Z(n860) );
  COND1XL U3000 ( .A(n3509), .B(n2322), .C(n2598), .Z(n858) );
  COND1XL U3001 ( .A(n3509), .B(n2321), .C(n2590), .Z(n866) );
  CANR2X1 U3002 ( .A(n3506), .B(n2418), .C(result[53]), .D(n3503), .Z(n2590)
         );
  COND1XL U3003 ( .A(n3510), .B(n4655), .C(n2591), .Z(n865) );
  CANR2X1 U3004 ( .A(n3506), .B(n4538), .C(result[54]), .D(n3503), .Z(n2591)
         );
  COND1XL U3005 ( .A(n3509), .B(n2316), .C(n2595), .Z(n861) );
  CANR2X1 U3006 ( .A(n3506), .B(n2335), .C(result[58]), .D(n3503), .Z(n2595)
         );
  COND1XL U3007 ( .A(n3509), .B(n2315), .C(n2545), .Z(n911) );
  CANR2X1 U3008 ( .A(n3507), .B(n2366), .C(result[8]), .D(n3504), .Z(n2545) );
  COND1XL U3009 ( .A(n3509), .B(n2314), .C(n2593), .Z(n863) );
  CANR2X1 U3010 ( .A(n3506), .B(n2334), .C(result[56]), .D(n3503), .Z(n2593)
         );
  COND1XL U3011 ( .A(n3510), .B(n2313), .C(n2581), .Z(n875) );
  COND1XL U3012 ( .A(n3510), .B(n2309), .C(n2559), .Z(n897) );
  COND1XL U3013 ( .A(n3509), .B(n3241), .C(n2553), .Z(n903) );
  CANR2X1 U3014 ( .A(n3507), .B(n2358), .C(result[16]), .D(n3505), .Z(n2553)
         );
  COND1XL U3015 ( .A(n3510), .B(n4143), .C(n2550), .Z(n906) );
  COND1XL U3016 ( .A(n3509), .B(n4154), .C(n2548), .Z(n908) );
  CANR2X1 U3017 ( .A(n3507), .B(n2364), .C(result[11]), .D(n3504), .Z(n2548)
         );
  COND1XL U3018 ( .A(n3509), .B(n4137), .C(n2544), .Z(n912) );
  CANR2X1 U3019 ( .A(n3507), .B(n2348), .C(result[7]), .D(n3504), .Z(n2544) );
  COND1XL U3020 ( .A(n3510), .B(n3203), .C(n2538), .Z(n918) );
  COND1XL U3021 ( .A(n3509), .B(n3264), .C(n2542), .Z(n914) );
  COND1XL U3022 ( .A(n3509), .B(n2369), .C(n3153), .Z(n793) );
  CANR2X1 U3023 ( .A(n3506), .B(n4660), .C(result[63]), .D(n3503), .Z(n3153)
         );
  COND1XL U3024 ( .A(n3407), .B(n3610), .C(n3609), .Z(n953) );
  CANR1XL U3025 ( .A(n4649), .B(n3608), .C(n3405), .Z(n3609) );
  COND1XL U3026 ( .A(n4661), .B(n3269), .C(n2439), .Z(n957) );
  CEOX1 U3027 ( .A(opera1[25]), .B(opera1[31]), .Z(n3427) );
  CND3X1 U3028 ( .A(n3518), .B(n3517), .C(n3516), .Z(n3522) );
  CND3X1 U3029 ( .A(n3374), .B(n3524), .C(n3523), .Z(n3528) );
  CEOX1 U3030 ( .A(opera1[21]), .B(n3512), .Z(n3428) );
  CEOX1 U3031 ( .A(opera1[22]), .B(n3215), .Z(n3429) );
  CND3XL U3032 ( .A(n3845), .B(n3844), .C(n3843), .Z(n840) );
  CANR1XL U3033 ( .A(result[48]), .B(n3200), .C(n3842), .Z(n3843) );
  CND2X1 U3034 ( .A(result[40]), .B(n3716), .Z(n3824) );
  CND3XL U3035 ( .A(n4129), .B(n4128), .C(n4127), .Z(n799) );
  CANR1XL U3036 ( .A(result[26]), .B(n3200), .C(n4126), .Z(n4127) );
  COND1XL U3037 ( .A(n4553), .B(n4012), .C(n4011), .Z(n831) );
  CNR2IX1 U3038 ( .B(result[58]), .A(n3501), .Z(n4008) );
  COND1XL U3039 ( .A(n3820), .B(n4553), .C(n3819), .Z(n833) );
  CEOX1 U3040 ( .A(opera1[23]), .B(opera1[31]), .Z(n3435) );
  CENX1 U3041 ( .A(opera1[26]), .B(n3353), .Z(n3437) );
  CND2X1 U3042 ( .A(valid), .B(n4394), .Z(n3583) );
  CAN2X1 U3043 ( .A(i[5]), .B(i[4]), .Z(n3438) );
  CND2XL U3044 ( .A(i[18]), .B(i[19]), .Z(n4606) );
  CND2X1 U3045 ( .A(res_not_wire[14]), .B(n1475), .Z(n4088) );
  CNR2IXL U3046 ( .B(result[36]), .A(n4495), .Z(n3601) );
  CND2X1 U3047 ( .A(result[61]), .B(n3401), .Z(n4058) );
  CND3XL U3048 ( .A(n3892), .B(n3891), .C(n3890), .Z(n855) );
  CANR1XL U3049 ( .A(result[33]), .B(n3200), .C(n3889), .Z(n3890) );
  CND3XL U3050 ( .A(n4465), .B(n4464), .C(n4463), .Z(n847) );
  CANR1XL U3051 ( .A(result[41]), .B(n3200), .C(n4462), .Z(n4463) );
  CND3XL U3052 ( .A(n4473), .B(n4472), .C(n4471), .Z(n846) );
  CANR1XL U3053 ( .A(result[42]), .B(n3200), .C(n4470), .Z(n4471) );
  CND3XL U3054 ( .A(n4111), .B(n4110), .C(n4109), .Z(n805) );
  CANR1XL U3055 ( .A(result[20]), .B(n3200), .C(n4108), .Z(n4109) );
  CND3XL U3056 ( .A(n3209), .B(n4333), .C(n4092), .Z(n4111) );
  CND3XL U3057 ( .A(n4375), .B(n4259), .C(n4136), .Z(n4142) );
  CANR1XL U3058 ( .A(result[8]), .B(n3200), .C(n4139), .Z(n4140) );
  CND3XL U3059 ( .A(n4159), .B(n4158), .C(n4157), .Z(n814) );
  CANR1XL U3060 ( .A(result[11]), .B(n3200), .C(n4156), .Z(n4157) );
  CND3XL U3061 ( .A(n4181), .B(n4180), .C(n4179), .Z(n819) );
  CND3XL U3062 ( .A(n4375), .B(n4175), .C(n4174), .Z(n4181) );
  CANR1XL U3063 ( .A(result[6]), .B(n3200), .C(n4178), .Z(n4179) );
  CND3XL U3064 ( .A(n4196), .B(n4195), .C(n4194), .Z(n813) );
  CANR1XL U3065 ( .A(result[12]), .B(n3200), .C(n4193), .Z(n4194) );
  CND3XL U3066 ( .A(n4248), .B(n4247), .C(n4246), .Z(n822) );
  CND3XL U3067 ( .A(n4245), .B(n4244), .C(n4375), .Z(n4246) );
  COND3XL U3068 ( .A(n1472), .B(n4240), .C(n4252), .D(n3211), .Z(n4247) );
  CANR2XL U3069 ( .A(result[4]), .B(n3500), .C(result[3]), .D(n3200), .Z(n4248) );
  CND3XL U3070 ( .A(n4268), .B(n4267), .C(n4266), .Z(n816) );
  CANR1XL U3071 ( .A(result[9]), .B(n3200), .C(n4265), .Z(n4266) );
  CND3XL U3072 ( .A(n4323), .B(n4322), .C(n4321), .Z(n810) );
  CANR1XL U3073 ( .A(result[15]), .B(n3200), .C(n4320), .Z(n4321) );
  CND3XL U3074 ( .A(n4382), .B(n4204), .C(n4375), .Z(n4205) );
  CANR1XL U3075 ( .A(result[29]), .B(n3200), .C(n4358), .Z(n4359) );
  CND3XL U3076 ( .A(n4087), .B(n4086), .C(n4085), .Z(n825) );
  CND2XL U3077 ( .A(n3211), .B(n4083), .Z(n4086) );
  CANR1XL U3078 ( .A(result[0]), .B(n3200), .C(n4084), .Z(n4085) );
  CND3XL U3079 ( .A(n4150), .B(n4149), .C(n4148), .Z(n811) );
  CND3XL U3080 ( .A(n3207), .B(n4318), .C(n4144), .Z(n4150) );
  CANR1XL U3081 ( .A(result[14]), .B(n3200), .C(n4147), .Z(n4148) );
  CND3XL U3082 ( .A(n4166), .B(n4165), .C(n4164), .Z(n823) );
  CND3XL U3083 ( .A(n3209), .B(n4167), .C(n4160), .Z(n4166) );
  CANR1XL U3084 ( .A(result[2]), .B(n3200), .C(n4163), .Z(n4164) );
  CND3XL U3085 ( .A(n4173), .B(n4172), .C(n4171), .Z(n821) );
  CND2XL U3086 ( .A(n3209), .B(n4168), .Z(n4173) );
  CANR1XL U3087 ( .A(result[4]), .B(n3200), .C(n4170), .Z(n4171) );
  CND3XL U3088 ( .A(n4187), .B(n4186), .C(n4185), .Z(n815) );
  CND2XL U3089 ( .A(n3209), .B(n4182), .Z(n4187) );
  CANR1XL U3090 ( .A(result[10]), .B(n3200), .C(n4184), .Z(n4185) );
  CND3XL U3091 ( .A(n4239), .B(n4238), .C(n4237), .Z(n824) );
  CND2XL U3092 ( .A(n3211), .B(n4232), .Z(n4239) );
  CND3XL U3093 ( .A(n4375), .B(n4243), .C(n4235), .Z(n4238) );
  CANR1XL U3094 ( .A(result[1]), .B(n3200), .C(n4236), .Z(n4237) );
  CND3XL U3095 ( .A(n4375), .B(n4251), .C(n4250), .Z(n4258) );
  CND3XL U3096 ( .A(n3209), .B(n4254), .C(n4253), .Z(n4257) );
  CANR1XL U3097 ( .A(result[5]), .B(n3200), .C(n4255), .Z(n4256) );
  CND3XL U3098 ( .A(n4277), .B(n4276), .C(n4275), .Z(n812) );
  CND2XL U3099 ( .A(n3211), .B(n4270), .Z(n4277) );
  CANR1XL U3100 ( .A(result[13]), .B(n3200), .C(n4274), .Z(n4275) );
  CND3XL U3101 ( .A(n4285), .B(n4284), .C(n4283), .Z(n818) );
  CND2XL U3102 ( .A(n3207), .B(n4279), .Z(n4285) );
  CANR1XL U3103 ( .A(result[7]), .B(n3200), .C(n4282), .Z(n4283) );
  CND3XL U3104 ( .A(n4332), .B(n4331), .C(n4330), .Z(n808) );
  CND3XL U3105 ( .A(n3211), .B(n4326), .C(n4325), .Z(n4332) );
  CANR1XL U3106 ( .A(result[17]), .B(n3200), .C(n4329), .Z(n4330) );
  CNR2IXL U3107 ( .B(result[58]), .A(n4495), .Z(n4413) );
  CNR2IXL U3108 ( .B(result[55]), .A(n4495), .Z(n3817) );
  CNR2IXL U3109 ( .B(result[61]), .A(n4495), .Z(n3795) );
  CND2IX1 U3110 ( .B(n114), .A(n3789), .Z(n3853) );
  CEOXL U3111 ( .A(opera2[10]), .B(n3195), .Z(n3443) );
  CND2X1 U3112 ( .A(n1128), .B(res_not_wire[52]), .Z(n3851) );
  CND2X1 U3113 ( .A(result[34]), .B(n3366), .Z(n4444) );
  CANR1XL U3114 ( .A(result[18]), .B(n3200), .C(n4219), .Z(n4220) );
  CND2X1 U3115 ( .A(res_not_wire[50]), .B(n3447), .Z(n3970) );
  CND2XL U3116 ( .A(result[32]), .B(n3200), .Z(n3920) );
  CANR1XL U3117 ( .A(n3603), .B(n3602), .C(n3601), .Z(n3604) );
  CNR2IXL U3118 ( .B(n4429), .A(n3509), .Z(n3895) );
  COND2XL U3119 ( .A(n3501), .B(n3221), .C(n4495), .D(n3244), .Z(n3905) );
  CNR2IXL U3120 ( .B(res_not_wire[36]), .A(n3509), .Z(n3907) );
  CANR2X1 U3121 ( .A(n3507), .B(n2359), .C(result[12]), .D(n3504), .Z(n2549)
         );
  CNR2IX1 U3122 ( .B(res_not_wire[12]), .A(n3510), .Z(n3934) );
  CNR2IX1 U3123 ( .B(n3226), .A(n3509), .Z(n3956) );
  CNR2IX1 U3124 ( .B(n3220), .A(n3510), .Z(n4072) );
  CNR2IX1 U3125 ( .B(res_not_wire[28]), .A(n3510), .Z(n4556) );
  CANR2X1 U3126 ( .A(n3508), .B(n2356), .C(result[28]), .D(n3413), .Z(n2565)
         );
  CNR2IX1 U3127 ( .B(res_not_wire[18]), .A(n3510), .Z(n4559) );
  CANR2X1 U3128 ( .A(n3507), .B(n2345), .C(result[15]), .D(n3504), .Z(n2552)
         );
  CNR2IX1 U3129 ( .B(n43), .A(n3510), .Z(n4560) );
  COND2XL U3130 ( .A(n3501), .B(n4474), .C(n4495), .D(n2329), .Z(n4486) );
  CND2X1 U3131 ( .A(n3448), .B(n3963), .Z(n887) );
  COR2XL U3132 ( .A(n3350), .B(n3509), .Z(n3448) );
  CND2X1 U3133 ( .A(n3449), .B(n4528), .Z(n885) );
  COR2XL U3134 ( .A(n2324), .B(n3509), .Z(n3449) );
  CNR2IX1 U3135 ( .B(n3254), .A(n3510), .Z(n3939) );
  CNR2IX1 U3136 ( .B(n3236), .A(n3510), .Z(n4543) );
  CANR2X1 U3137 ( .A(n3507), .B(n2350), .C(result[9]), .D(n3504), .Z(n2546) );
  CNR2IX1 U3138 ( .B(n1474), .A(n3509), .Z(n3935) );
  CMXI2X1 U3139 ( .A0(n3959), .A1(n3960), .S(i[3]), .Z(n3961) );
  CNR2IXL U3140 ( .B(n1472), .A(n3510), .Z(n3962) );
  CND2XL U3141 ( .A(i[15]), .B(i[28]), .Z(n3576) );
  CND2X1 U3142 ( .A(n43), .B(n4343), .Z(n3594) );
  CND2XL U3143 ( .A(i[20]), .B(i[21]), .Z(n3573) );
  CND2X1 U3144 ( .A(res_not_wire[28]), .B(n4356), .Z(n3593) );
  CEOX2 U3145 ( .A(opera1[12]), .B(opera1[31]), .Z(n3451) );
  CIVX2 U3146 ( .A(n3587), .Z(n4176) );
  CND2X1 U3147 ( .A(n3445), .B(n3958), .Z(n3960) );
  CENX1 U3148 ( .A(opera1[29]), .B(opera1[31]), .Z(n3628) );
  CENX1 U3149 ( .A(res_not_wire[10]), .B(n4264), .Z(n4182) );
  CENX1 U3150 ( .A(opera2[22]), .B(n3197), .Z(n4115) );
  COND1XL U3151 ( .A(n4252), .B(n3225), .C(n2382), .Z(n4253) );
  CND2XL U3152 ( .A(n1472), .B(n4240), .Z(n4252) );
  CNR2IXL U3153 ( .B(i[24]), .A(n4624), .Z(n4626) );
  CND2XL U3154 ( .A(res_not_wire[38]), .B(n3821), .Z(n3941) );
  CEOXL U3155 ( .A(c_inres), .B(res_not_wire[0]), .Z(n4083) );
  CNR2X1 U3156 ( .A(n3288), .B(nst[0]), .Z(n55) );
  CNR2X1 U3157 ( .A(n3288), .B(n2336), .Z(N34) );
  CND2XL U3158 ( .A(n3655), .B(n3654), .Z(n3656) );
  COND1X1 U3159 ( .A(n3720), .B(n3293), .C(n3719), .Z(n3722) );
  CIVXL U3160 ( .A(n3719), .Z(n3715) );
  CIVX1 U3161 ( .A(n3964), .Z(n3967) );
  CANR2XL U3162 ( .A(result[25]), .B(n3500), .C(result[24]), .D(n3200), .Z(
        n4207) );
  CNR2IXL U3163 ( .B(n4402), .A(n4396), .Z(n4408) );
  CIVX1 U3164 ( .A(n4396), .Z(n4005) );
  CND2IX1 U3165 ( .B(n3416), .A(n3768), .Z(n3690) );
  CENX1 U3166 ( .A(n3995), .B(n3994), .Z(n4001) );
  COND1X2 U3167 ( .A(n3778), .B(n3808), .C(n3216), .Z(n3779) );
  CIVX2 U3168 ( .A(n3689), .Z(n4491) );
  CIVXL U3169 ( .A(n4054), .Z(n4055) );
  CENX1 U3170 ( .A(n3786), .B(n4015), .Z(n4020) );
  CIVXL U3171 ( .A(n3430), .Z(n3468) );
  CANR1XL U3172 ( .A(n3315), .B(n3455), .C(n3457), .Z(n4216) );
  CANR1XL U3173 ( .A(n3396), .B(n4439), .C(n4429), .Z(n4438) );
  CND2X1 U3174 ( .A(n4221), .B(n4220), .Z(n807) );
  CMXI2XL U3175 ( .A0(n4635), .A1(n4634), .S(i[26]), .Z(n928) );
  CANR11XL U3176 ( .A(n3207), .B(n4370), .C(n4218), .D(n4217), .Z(n4221) );
  CND2XL U3177 ( .A(i[26]), .B(i[27]), .Z(n4641) );
  CND2X1 U3178 ( .A(n3520), .B(n3519), .Z(n3521) );
  CEOXL U3179 ( .A(opera1[6]), .B(n3512), .Z(n3471) );
  CNIVX1 U3180 ( .A(n3848), .Z(n3472) );
  CND2XL U3181 ( .A(n4421), .B(n3480), .Z(n3473) );
  CANR1X2 U3182 ( .A(n3738), .B(n3825), .C(n3802), .Z(n3740) );
  CND2XL U3183 ( .A(n3367), .B(n3713), .Z(n3719) );
  CND2XL U3184 ( .A(n4152), .B(n4151), .Z(n4153) );
  CNR2X1 U3185 ( .A(n4028), .B(n4027), .Z(n4029) );
  CND2IXL U3186 ( .B(n4529), .A(n4419), .Z(n3489) );
  CND3XL U3187 ( .A(n4312), .B(n4311), .C(n4310), .Z(n802) );
  CND3XL U3188 ( .A(n3211), .B(n4269), .C(n4192), .Z(n4195) );
  CND3XL U3189 ( .A(n3211), .B(n4191), .C(n4155), .Z(n4158) );
  COND1XL U3190 ( .A(n4269), .B(n4143), .C(n3247), .Z(n4144) );
  CIVX1 U3191 ( .A(n4294), .Z(n4293) );
  CND2X1 U3192 ( .A(n3561), .B(n3618), .Z(n3562) );
  CND2XL U3193 ( .A(n3502), .B(n4293), .Z(n4296) );
  CENXL U3194 ( .A(n3193), .B(n3215), .Z(n3612) );
  CND2XL U3195 ( .A(n3640), .B(n3639), .Z(n3764) );
  CIVX1 U3196 ( .A(n3764), .Z(n3641) );
  CND2X2 U3197 ( .A(n3710), .B(n3478), .Z(n3698) );
  CNIVXL U3198 ( .A(n3486), .Z(n3478) );
  COND1XL U3199 ( .A(n4639), .B(n4645), .C(n4638), .Z(n927) );
  COND1XL U3200 ( .A(n4598), .B(n4645), .C(n4597), .Z(n939) );
  COND1XL U3201 ( .A(n4568), .B(n4645), .C(n4567), .Z(n947) );
  CMXI2XL U3202 ( .A0(n4645), .A1(n4642), .S(i[0]), .Z(n952) );
  COND2XL U3203 ( .A(n4642), .B(n4513), .C(n4512), .D(n4645), .Z(n955) );
  CAOR2XL U3204 ( .A(n3509), .B(n4653), .C(valid), .D(n3217), .Z(n923) );
  CND2XL U3205 ( .A(n4623), .B(n4622), .Z(n4627) );
  CND2XL U3206 ( .A(n4623), .B(n4610), .Z(n4611) );
  COND1XL U3207 ( .A(n4633), .B(n4645), .C(n4642), .Z(n4637) );
  COND1XL U3208 ( .A(n4615), .B(n4645), .C(n4642), .Z(n4618) );
  COND1XL U3209 ( .A(n4593), .B(n4645), .C(n4642), .Z(n4596) );
  COND1XL U3210 ( .A(n4563), .B(n4645), .C(n4642), .Z(n4566) );
  COND1XL U3211 ( .A(n4645), .B(i[17]), .C(n3454), .Z(n4603) );
  CND3XL U3212 ( .A(result[0]), .B(n4653), .C(n3232), .Z(n3918) );
  CND3XL U3213 ( .A(n53), .B(n2060), .C(n3513), .Z(n4661) );
  CND3XL U3214 ( .A(n4375), .B(n3314), .C(n4198), .Z(n4201) );
  CND2XL U3215 ( .A(n4272), .B(n4271), .Z(n4273) );
  CENX1 U3216 ( .A(result[57]), .B(n3761), .Z(n3480) );
  CENX1 U3217 ( .A(opera1[20]), .B(n3215), .Z(n3652) );
  CND4X2 U3218 ( .A(n3352), .B(n3492), .C(n3486), .D(n3493), .Z(n3619) );
  CANR1X1 U3219 ( .A(n4069), .B(n4070), .C(n4068), .Z(n4659) );
  CND3XL U3220 ( .A(n3211), .B(n4264), .C(n4263), .Z(n4267) );
  CND3XL U3221 ( .A(n3211), .B(n4365), .C(n4364), .Z(n4368) );
  COND1XL U3222 ( .A(n4264), .B(n3253), .C(n4154), .Z(n4155) );
  CND2XL U3223 ( .A(n4065), .B(n4417), .Z(n4396) );
  CND2XL U3224 ( .A(n4042), .B(n4417), .Z(n4399) );
  CENX1 U3225 ( .A(result[57]), .B(n3761), .Z(n3485) );
  CANR1XL U3226 ( .A(n3636), .B(n3638), .C(n3324), .Z(n3481) );
  CND2IX2 U3227 ( .B(n3864), .A(n3325), .Z(n3898) );
  COND3X1 U3228 ( .A(n3858), .B(n4553), .C(n3857), .D(n3856), .Z(n835) );
  COND3X1 U3229 ( .A(n3933), .B(n4553), .C(n3932), .D(n3931), .Z(n843) );
  CND2IX1 U3230 ( .B(n3990), .A(n3980), .Z(n3759) );
  CND2IX2 U3231 ( .B(n4028), .A(n3979), .Z(n3483) );
  CND3XL U3232 ( .A(n4375), .B(n4234), .C(n4082), .Z(n4087) );
  CND2XL U3233 ( .A(n4234), .B(n4233), .Z(n4235) );
  CND2IXL U3234 ( .B(c_inop2), .A(n4081), .Z(n4082) );
  CND2XL U3235 ( .A(n4372), .B(n4371), .Z(n4373) );
  COND3XL U3236 ( .A(n4391), .B(n2337), .C(n4661), .D(n4390), .Z(n922) );
  COND4CXL U3237 ( .A(n4420), .B(n4419), .C(n4418), .D(n4417), .Z(n4421) );
  COND3X1 U3238 ( .A(n4541), .B(n4553), .C(n4540), .D(n4539), .Z(n834) );
  CND2XL U3239 ( .A(n3867), .B(n3924), .Z(n3926) );
  CND3XL U3240 ( .A(n3211), .B(n4262), .C(n4138), .Z(n4141) );
  COND3X1 U3241 ( .A(n4122), .B(res_not_wire[24]), .C(n4380), .D(n3207), .Z(
        n4206) );
  CND2IXL U3242 ( .B(n1474), .A(n4262), .Z(n4263) );
  CND3XL U3243 ( .A(c_inres), .B(n3218), .C(n4176), .Z(n4254) );
  CND3X1 U3244 ( .A(res_not_wire[20]), .B(n4223), .C(n3230), .Z(n4333) );
  CND2XL U3245 ( .A(c_inres), .B(res_not_wire[0]), .Z(n4231) );
  COND3X1 U3246 ( .A(n4428), .B(n4553), .C(n4427), .D(n4426), .Z(n832) );
  CND2IX2 U3247 ( .B(n3846), .A(n3780), .Z(n4419) );
  CND2X1 U3248 ( .A(n3985), .B(n4402), .Z(n3757) );
  CND2X1 U3249 ( .A(n3481), .B(result[56]), .Z(n4417) );
  CND2XL U3250 ( .A(n3363), .B(n4019), .Z(n4022) );
  CND2X1 U3251 ( .A(n3751), .B(n3745), .Z(n3746) );
  CND2IX2 U3252 ( .B(n3809), .A(n3966), .Z(n3808) );
  CND3XL U3253 ( .A(n4375), .B(n4353), .C(n4346), .Z(n4349) );
  CND3XL U3254 ( .A(n4375), .B(n4374), .C(n4373), .Z(n4378) );
  COND1XL U3255 ( .A(n4353), .B(n4352), .C(n3272), .Z(n4354) );
  COND1XL U3256 ( .A(n4374), .B(n4336), .C(n4335), .Z(n4337) );
  CNR2XL U3257 ( .A(n4130), .B(n4242), .Z(n4131) );
  CND2X1 U3258 ( .A(n3363), .B(n4417), .Z(n3763) );
  CIVDX1 U3259 ( .A(n3652), .Z0(n3488), .Z1(n3487) );
  CANR1XL U3260 ( .A(n3441), .B(n3944), .C(n3945), .Z(n3908) );
  CND3XL U3261 ( .A(n3209), .B(n3377), .C(n4177), .Z(n4180) );
  COND1XL U3262 ( .A(n3377), .B(n4137), .C(n3248), .Z(n4138) );
  CNR2IXL U3263 ( .B(n4363), .A(n3208), .Z(n4355) );
  CND2XL U3264 ( .A(n4481), .B(n3447), .Z(n3972) );
  CND2XL U3265 ( .A(n4481), .B(n3871), .Z(n4469) );
  CND2IX2 U3266 ( .B(n4529), .A(n4419), .Z(n4044) );
  CND2IXL U3267 ( .B(n3452), .A(n3566), .Z(n3564) );
  CND3XL U3268 ( .A(n3367), .B(n3303), .C(n3633), .Z(n3490) );
  CIVXL U3269 ( .A(n3556), .Z(n3561) );
  CND3XL U3270 ( .A(n4375), .B(n3312), .C(n4273), .Z(n4276) );
  CND3XL U3271 ( .A(n4375), .B(n4362), .C(n4354), .Z(n4361) );
  COND1XL U3272 ( .A(n4315), .B(n3312), .C(n4313), .Z(n4316) );
  CND4XL U3273 ( .A(n4133), .B(n4132), .C(n4131), .D(n4161), .Z(n4259) );
  CNR2XL U3274 ( .A(n3683), .B(n3682), .Z(n3686) );
  CND2X1 U3275 ( .A(n3367), .B(n3718), .Z(n3730) );
  CND2IXL U3276 ( .B(result[55]), .A(n3706), .Z(n3707) );
  CIVX1 U3277 ( .A(n4042), .Z(n4025) );
  CND3X1 U3278 ( .A(n3701), .B(n3675), .C(n3368), .Z(n3700) );
  COND3X1 U3279 ( .A(n4511), .B(n4553), .C(n4510), .D(n4509), .Z(n837) );
  CIVXL U3280 ( .A(n3294), .Z(n4400) );
  COND1X1 U3281 ( .A(n3661), .B(n3451), .C(n3669), .Z(n3693) );
  CND3XL U3282 ( .A(n3211), .B(n4324), .C(n4319), .Z(n4322) );
  COND3XL U3283 ( .A(n4305), .B(n4304), .C(n3207), .D(n4303), .Z(n4312) );
  COND1XL U3284 ( .A(n4324), .B(n3241), .C(n148), .Z(n4325) );
  CNR3XL U3285 ( .A(n4324), .B(n4209), .C(n138), .Z(n4357) );
  CND2X1 U3286 ( .A(n3472), .B(n3847), .Z(n3878) );
  CND2IX2 U3287 ( .B(n4457), .A(n3726), .Z(n3802) );
  CND2XL U3288 ( .A(n3755), .B(n3749), .Z(n3750) );
  CND2X1 U3289 ( .A(n3642), .B(n3644), .Z(n3771) );
  CIVX1 U3290 ( .A(n4397), .Z(n4406) );
  CIVDX2 U3291 ( .A(n3657), .Z0(n3495), .Z1(n3494) );
  CNR3X2 U3292 ( .A(n3632), .B(n3654), .C(n3631), .Z(n3633) );
  CND2X1 U3293 ( .A(n3687), .B(n3688), .Z(n3769) );
  COND1X1 U3294 ( .A(n3712), .B(n3478), .C(n3711), .Z(n3723) );
  CND2X1 U3295 ( .A(result[37]), .B(n3728), .Z(n3732) );
  CND2IXL U3296 ( .B(n3429), .A(n3648), .Z(n3639) );
  CND2IXL U3297 ( .B(n3428), .A(n3490), .Z(n3647) );
  CND2IXL U3298 ( .B(n3435), .A(n3640), .Z(n3637) );
  COND3X1 U3299 ( .A(n4039), .B(n4553), .C(n4038), .D(n4037), .Z(n826) );
  COND3X1 U3300 ( .A(n4301), .B(n4384), .C(n4300), .D(n4299), .Z(n794) );
  CND3XL U3301 ( .A(n4375), .B(n4189), .C(n4153), .Z(n4159) );
  CND3XL U3302 ( .A(n4375), .B(n4317), .C(n4316), .Z(n4323) );
  CND3XL U3303 ( .A(n4375), .B(n3327), .C(n4260), .Z(n4268) );
  CND2XL U3304 ( .A(n4189), .B(n4188), .Z(n4190) );
  CND2XL U3305 ( .A(n4317), .B(n4197), .Z(n4198) );
  CNR3XL U3306 ( .A(n4216), .B(n4215), .C(n4384), .Z(n4217) );
  CND2X1 U3307 ( .A(n4003), .B(n3295), .Z(n4418) );
  CANR1XL U3308 ( .A(n4025), .B(n3430), .C(n4028), .Z(n4026) );
  COND3X1 U3309 ( .A(n4403), .B(n3294), .C(n4401), .D(n4402), .Z(n4405) );
  CIVXL U3310 ( .A(n3500), .Z(n3499) );
  CIVX2 U3311 ( .A(n3291), .Z(n4654) );
  CIVX2 U3312 ( .A(n4661), .Z(n4079) );
  CIVX2 U3313 ( .A(n3514), .Z(n3584) );
  CIVX2 U3314 ( .A(n3543), .Z(n4653) );
  CIVX2 U3315 ( .A(i[22]), .Z(n3518) );
  CNR3X2 U3316 ( .A(i[28]), .B(i[30]), .C(i[29]), .Z(n3520) );
  CNR3X2 U3317 ( .A(i[25]), .B(i[27]), .C(i[26]), .Z(n3519) );
  CNR3X2 U3318 ( .A(i[15]), .B(i[18]), .C(i[17]), .Z(n3526) );
  CNR3X2 U3319 ( .A(i[12]), .B(i[14]), .C(i[13]), .Z(n3525) );
  CNR2X2 U3320 ( .A(n3527), .B(n3528), .Z(n3529) );
  CND2X2 U3321 ( .A(n3530), .B(n3529), .Z(n3531) );
  CIVX2 U3322 ( .A(n3531), .Z(n3537) );
  CIVX2 U3323 ( .A(n3535), .Z(n3544) );
  CIVX2 U3324 ( .A(i[16]), .Z(n3538) );
  CIVX2 U3325 ( .A(i[5]), .Z(n3610) );
  CND4X2 U3326 ( .A(n3538), .B(n3537), .C(n3610), .D(n3536), .Z(n3539) );
  CIVX2 U3327 ( .A(n3542), .Z(n3540) );
  CIVX2 U3328 ( .A(result[63]), .Z(n4660) );
  CIVX2 U3329 ( .A(n1476), .Z(n2369) );
  CIVX2 U3330 ( .A(res_not_wire[60]), .Z(n4657) );
  CIVX2 U3331 ( .A(result[59]), .Z(n2380) );
  CIVX2 U3332 ( .A(result[58]), .Z(n2335) );
  CIVX2 U3333 ( .A(res_not_wire[54]), .Z(n4655) );
  CIVX2 U3334 ( .A(res_not_wire[48]), .Z(n4658) );
  CIVX2 U3335 ( .A(result[31]), .Z(n2347) );
  CIVX2 U3336 ( .A(result[0]), .Z(n4656) );
  CND2IX1 U3337 ( .B(n3543), .A(n3542), .Z(n4390) );
  CND2IX1 U3338 ( .B(n3544), .A(n4390), .Z(n3549) );
  CIVX2 U3339 ( .A(n4391), .Z(n4393) );
  CMXI2X1 U3340 ( .A0(n4394), .A1(nst[0]), .S(n4393), .Z(n2439) );
  CIVX2 U3341 ( .A(n3549), .Z(n3550) );
  CIVX2 U3342 ( .A(n4569), .Z(n4571) );
  CIVX2 U3343 ( .A(n4588), .Z(n4582) );
  CIVX2 U3344 ( .A(n4594), .Z(n4593) );
  CIVX2 U3345 ( .A(n3552), .Z(n4631) );
  CIVX2 U3346 ( .A(n3729), .Z(n3553) );
  CIVX2 U3347 ( .A(n3555), .Z(n3559) );
  CIVX2 U3348 ( .A(n3562), .Z(n3560) );
  CIVX2 U3349 ( .A(n4431), .Z(n3572) );
  CIVX2 U3350 ( .A(n4444), .Z(n3571) );
  CIVX2 U3351 ( .A(n3887), .Z(n4443) );
  CND2X2 U3352 ( .A(n3572), .B(n4432), .Z(n3727) );
  CIVX2 U3353 ( .A(n4390), .Z(n3581) );
  CIVX2 U3354 ( .A(n4624), .Z(n4632) );
  COND2X1 U3355 ( .A(n3582), .B(n4553), .C(n3501), .D(n3442), .Z(n3605) );
  CIVX2 U3356 ( .A(n130), .Z(n4429) );
  CND2IX1 U3357 ( .B(n3240), .A(n3585), .Z(n3586) );
  CIVX2 U3358 ( .A(n3586), .Z(n3821) );
  CIVX2 U3359 ( .A(n4278), .Z(n3588) );
  CIVX2 U3360 ( .A(n4191), .Z(n4089) );
  CIVX2 U3361 ( .A(n148), .Z(n4090) );
  CIVX2 U3362 ( .A(n142), .Z(n4304) );
  CIVX2 U3363 ( .A(n144), .Z(n4334) );
  CIVX2 U3364 ( .A(n3592), .Z(n4123) );
  CIVX2 U3365 ( .A(n4209), .Z(n3597) );
  CIVX2 U3366 ( .A(n136), .Z(n4356) );
  CIVX2 U3367 ( .A(n138), .Z(n4343) );
  CIVX2 U3368 ( .A(n3600), .Z(n4439) );
  CND2IX1 U3369 ( .B(n3606), .A(n2543), .Z(n913) );
  CND2IX1 U3370 ( .B(n3613), .A(n2563), .Z(n893) );
  CIVX2 U3371 ( .A(n3670), .Z(n3614) );
  CIVX2 U3372 ( .A(n3619), .Z(n3665) );
  CND2X2 U3373 ( .A(n3660), .B(n3416), .Z(n3620) );
  CIVX2 U3374 ( .A(n3620), .Z(n3634) );
  CIVX2 U3375 ( .A(n3654), .Z(n3622) );
  CIVX2 U3376 ( .A(n3636), .Z(n3635) );
  CIVX2 U3377 ( .A(n3749), .Z(n3623) );
  CIVX2 U3378 ( .A(n3751), .Z(n3626) );
  CIVX2 U3379 ( .A(n3745), .Z(n3625) );
  CND2X2 U3380 ( .A(n3626), .B(n3625), .Z(n3747) );
  CIVX2 U3381 ( .A(n3628), .Z(n3627) );
  CIVX2 U3382 ( .A(n3744), .Z(n3629) );
  CIVX2 U3383 ( .A(n3763), .Z(n3762) );
  CND2X2 U3384 ( .A(result[54]), .B(n3641), .Z(n3988) );
  CND2X2 U3385 ( .A(n3495), .B(n3415), .Z(n3644) );
  CND2X2 U3386 ( .A(n3645), .B(n3397), .Z(n3651) );
  CIVX2 U3387 ( .A(n3653), .Z(n3810) );
  CIVX2 U3388 ( .A(n3700), .Z(n3661) );
  CIVX2 U3389 ( .A(n3693), .Z(n3662) );
  CND2X2 U3390 ( .A(n3662), .B(result[44]), .Z(n3859) );
  CIVX2 U3391 ( .A(n3681), .Z(n3672) );
  CND2X2 U3392 ( .A(n3672), .B(result[45]), .Z(n3924) );
  CND2X2 U3393 ( .A(n3859), .B(n3924), .Z(n4477) );
  CIVX2 U3394 ( .A(n3680), .Z(n3927) );
  CIVX2 U3395 ( .A(n3804), .Z(n3691) );
  CIVX2 U3396 ( .A(n3696), .Z(n3713) );
  CND2X2 U3397 ( .A(n3479), .B(n3713), .Z(n3697) );
  CND2X2 U3398 ( .A(n4042), .B(n3707), .Z(n3811) );
  CIVX2 U3399 ( .A(n3711), .Z(n3709) );
  CIVX2 U3400 ( .A(n3803), .Z(n3738) );
  CIVX2 U3401 ( .A(n3717), .Z(n4520) );
  CIVX2 U3402 ( .A(n3730), .Z(n3720) );
  CENX2 U3403 ( .A(result[42]), .B(n3323), .Z(n4457) );
  CIVX2 U3404 ( .A(n3725), .Z(n4458) );
  CIVX2 U3405 ( .A(n3727), .Z(n3731) );
  CIVX2 U3406 ( .A(n3732), .Z(n3945) );
  COND1X2 U3407 ( .A(n3945), .B(n3441), .C(n3348), .Z(n3734) );
  CIVX2 U3408 ( .A(n3734), .Z(n3943) );
  CIVX2 U3409 ( .A(n3734), .Z(n3736) );
  CND2X2 U3410 ( .A(n3740), .B(n3739), .Z(n3861) );
  CND2X2 U3411 ( .A(n3743), .B(n3742), .Z(n4403) );
  CND2X2 U3412 ( .A(n4403), .B(n4042), .Z(n4003) );
  CIVX2 U3413 ( .A(n3985), .Z(n3990) );
  CIVX2 U3414 ( .A(n3760), .Z(n3756) );
  CIVX2 U3415 ( .A(n3981), .Z(n4007) );
  CIVX2 U3416 ( .A(n4027), .Z(n4420) );
  CND2IX1 U3417 ( .B(result[51]), .A(n3214), .Z(n3765) );
  CIVX2 U3418 ( .A(n3472), .Z(n3778) );
  COND4CX1 U3419 ( .A(n3472), .B(n3806), .C(n3779), .D(n3849), .Z(n3780) );
  CIVX2 U3420 ( .A(n4013), .Z(n4016) );
  CENX1 U3421 ( .A(result[62]), .B(n4016), .Z(n3786) );
  CIVX2 U3422 ( .A(n128), .Z(n3940) );
  CANR3X1 U3423 ( .A(n3209), .B(n3796), .C(n3795), .D(n3794), .Z(n3797) );
  CND2X2 U3424 ( .A(n3799), .B(n3800), .Z(n3823) );
  CND2X2 U3425 ( .A(n3801), .B(n3823), .Z(n3832) );
  CIVX2 U3426 ( .A(n3811), .Z(n4533) );
  CANR3X1 U3427 ( .A(n3209), .B(n3818), .C(n3817), .D(n3816), .Z(n3819) );
  CND2IX1 U3428 ( .B(n4553), .A(n3826), .Z(n3829) );
  COND3X1 U3429 ( .A(n3830), .B(n3210), .C(n3829), .D(n3828), .Z(n848) );
  COND3X1 U3430 ( .A(n3408), .B(res_not_wire[48]), .C(n3211), .D(n3972), .Z(
        n3844) );
  CIVX2 U3431 ( .A(n3859), .Z(n3865) );
  CND2X2 U3432 ( .A(n3861), .B(n3860), .Z(n4467) );
  CIVX2 U3433 ( .A(n4467), .Z(n3863) );
  CND2IX1 U3434 ( .B(n3865), .A(n3898), .Z(n3866) );
  CIVX2 U3435 ( .A(n3866), .Z(n3925) );
  CIVX2 U3436 ( .A(n3870), .Z(n3928) );
  CIVX2 U3437 ( .A(n4469), .Z(n3900) );
  CND2X1 U3438 ( .A(n3873), .B(n3872), .Z(n3876) );
  CND2IX1 U3439 ( .B(n3208), .A(n3880), .Z(n3883) );
  CEN3X2 U3440 ( .A(result[34]), .B(n3366), .C(n3887), .Z(n3888) );
  CMXI2X1 U3441 ( .A0(n3508), .A1(n3505), .S(result[40]), .Z(n3893) );
  CND2IX1 U3442 ( .B(n3895), .A(n3894), .Z(n884) );
  CND2IX1 U3443 ( .B(n3897), .A(n3896), .Z(n877) );
  CIVX2 U3444 ( .A(n3898), .Z(n4478) );
  CENX1 U3445 ( .A(n122), .B(n3900), .Z(n3901) );
  CANR2X1 U3446 ( .A(n3903), .B(n3902), .C(n3211), .D(n3901), .Z(n3904) );
  CND2IX1 U3447 ( .B(n3905), .A(n3904), .Z(n845) );
  CND2IX1 U3448 ( .B(n3907), .A(n3906), .Z(n883) );
  CENX1 U3449 ( .A(n3402), .B(n3940), .Z(n3913) );
  CND2IX1 U3450 ( .B(n4553), .A(n3909), .Z(n3912) );
  CENX1 U3451 ( .A(n3968), .B(n3350), .Z(n3923) );
  CMXI2X1 U3452 ( .A0(n3918), .A1(n3917), .S(n3916), .Z(n3919) );
  COND3X1 U3453 ( .A(n3923), .B(n3496), .C(n3922), .D(n3921), .Z(n856) );
  CENX1 U3454 ( .A(n120), .B(n3928), .Z(n3929) );
  CND2IX1 U3455 ( .B(n3394), .A(n3929), .Z(n3932) );
  CND2IX1 U3456 ( .B(n3934), .A(n2549), .Z(n907) );
  CND2IX1 U3457 ( .B(n3935), .A(n2546), .Z(n910) );
  CMXI2X1 U3458 ( .A0(n3508), .A1(n3505), .S(result[38]), .Z(n3936) );
  CMXI2X1 U3459 ( .A0(n3508), .A1(n3505), .S(result[50]), .Z(n3937) );
  CND2IX1 U3460 ( .B(n3939), .A(n3938), .Z(n872) );
  CIVX2 U3461 ( .A(n3942), .Z(n4517) );
  CENX1 U3462 ( .A(n4517), .B(n3948), .Z(n3949) );
  CND2IX1 U3463 ( .B(n4553), .A(n3949), .Z(n3952) );
  COND3X1 U3464 ( .A(n3954), .B(n3953), .C(n3952), .D(n3951), .Z(n850) );
  CND2IX1 U3465 ( .B(n3956), .A(n3955), .Z(n870) );
  CND2IX1 U3466 ( .B(i[2]), .A(n4649), .Z(n3958) );
  CND2IX1 U3467 ( .B(n3405), .A(n3961), .Z(n954) );
  CND2IX1 U3468 ( .B(n3962), .A(n2540), .Z(n916) );
  CMXI2X1 U3469 ( .A0(n3508), .A1(n3505), .S(result[32]), .Z(n3963) );
  CENX1 U3470 ( .A(n4504), .B(n3322), .Z(n3978) );
  CIVX2 U3471 ( .A(n3971), .Z(n4506) );
  CIVX2 U3472 ( .A(n3972), .Z(n4548) );
  CND2X1 U3473 ( .A(n3974), .B(n3973), .Z(n3977) );
  CIVX2 U3474 ( .A(n3982), .Z(n3983) );
  CIVX2 U3475 ( .A(n4417), .Z(n4028) );
  CIVX2 U3476 ( .A(n3988), .Z(n4529) );
  CIVX2 U3477 ( .A(n4065), .Z(n4398) );
  CIVX2 U3478 ( .A(result[62]), .Z(n4014) );
  CIVX2 U3479 ( .A(n4018), .Z(n4021) );
  CIVX2 U3480 ( .A(n3489), .Z(n4050) );
  CIVX2 U3481 ( .A(n4404), .Z(n4062) );
  CND2IX1 U3482 ( .B(n4072), .A(n4071), .Z(n876) );
  CMXI2X1 U3483 ( .A0(n3508), .A1(n3505), .S(result[52]), .Z(n4073) );
  CND2IX1 U3484 ( .B(n4078), .A(n4077), .Z(n878) );
  CIVX2 U3485 ( .A(n4081), .Z(n4080) );
  CIVX2 U3486 ( .A(res_not_wire[20]), .Z(n4091) );
  CIVX2 U3487 ( .A(n4234), .Z(n4094) );
  CIVX2 U3488 ( .A(n4233), .Z(n4093) );
  CIVX2 U3489 ( .A(n4243), .Z(n4161) );
  CIVX2 U3490 ( .A(n4280), .Z(n4097) );
  CND3X2 U3491 ( .A(n3199), .B(n3328), .C(n3440), .Z(n4130) );
  CIVX2 U3492 ( .A(n4261), .Z(n4098) );
  CIVX2 U3493 ( .A(n4151), .Z(n4099) );
  CIVX2 U3494 ( .A(n4188), .Z(n4100) );
  CIVX2 U3495 ( .A(n4272), .Z(n4103) );
  CIVX2 U3496 ( .A(n4271), .Z(n4102) );
  CND2X2 U3497 ( .A(n4103), .B(n4102), .Z(n4314) );
  CIVX2 U3498 ( .A(n4313), .Z(n4104) );
  CIVX2 U3499 ( .A(n4315), .Z(n4145) );
  CIVX2 U3500 ( .A(n4197), .Z(n4105) );
  CIVX2 U3501 ( .A(n4372), .Z(n4215) );
  CIVX2 U3502 ( .A(n4371), .Z(n4106) );
  CND2X2 U3503 ( .A(n4215), .B(n4106), .Z(n4374) );
  CND2IX1 U3504 ( .B(n4384), .A(n4107), .Z(n4110) );
  CIVX2 U3505 ( .A(n4335), .Z(n4117) );
  CIVX2 U3506 ( .A(n4336), .Z(n4116) );
  CIVX2 U3507 ( .A(n4303), .Z(n4122) );
  CIVX2 U3508 ( .A(n4380), .Z(n4125) );
  COND4CX1 U3509 ( .A(n38), .B(n4125), .C(res_not_wire[26]), .D(n4124), .Z(
        n4128) );
  CIVX2 U3510 ( .A(n4134), .Z(n4132) );
  CIVX2 U3511 ( .A(n1891), .Z(n4137) );
  CIVX2 U3512 ( .A(n1475), .Z(n4143) );
  CIVX2 U3513 ( .A(n1918), .Z(n4154) );
  CIVX2 U3514 ( .A(n4167), .Z(n4240) );
  CND2IX1 U3515 ( .B(n3199), .A(n4251), .Z(n4174) );
  CIVX2 U3516 ( .A(n4344), .Z(n4208) );
  CND2IX1 U3517 ( .B(n3212), .A(n4210), .Z(n4213) );
  COND3X1 U3518 ( .A(n4230), .B(n3496), .C(n4229), .D(n4228), .Z(n803) );
  CENX1 U3519 ( .A(n1849), .B(n4231), .Z(n4232) );
  CND2IX1 U3520 ( .B(n3417), .A(n4259), .Z(n4260) );
  CIVX2 U3521 ( .A(n4351), .Z(n4287) );
  CENX1 U3522 ( .A(n134), .B(n4291), .Z(n4292) );
  CND2X1 U3523 ( .A(n3211), .B(n4292), .Z(n4300) );
  CND2IX1 U3524 ( .B(n2347), .A(n3200), .Z(n4298) );
  CMXI2X1 U3525 ( .A0(n4296), .A1(n4295), .S(result[32]), .Z(n4297) );
  CENX1 U3526 ( .A(n3404), .B(n4343), .Z(n4350) );
  COND4CX1 U3527 ( .A(res_not_wire[28]), .B(n4357), .C(n4356), .D(n4355), .Z(
        n4360) );
  COND3X1 U3528 ( .A(n4369), .B(n4384), .C(n4368), .D(n4367), .Z(n795) );
  CENX1 U3529 ( .A(n146), .B(n4370), .Z(n4379) );
  CENX1 U3530 ( .A(n4380), .B(n3229), .Z(n4389) );
  COND3X1 U3531 ( .A(n4389), .B(n3212), .C(n4388), .D(n4387), .Z(n800) );
  CMXI2X1 U3532 ( .A0(n4394), .A1(nst[2]), .S(n4393), .Z(n4395) );
  CANR3X1 U3533 ( .A(n3209), .B(n4414), .C(n4413), .D(n4412), .Z(n4415) );
  CND2IX1 U3534 ( .B(n2334), .A(n3200), .Z(n4426) );
  CND2IX1 U3535 ( .B(n3394), .A(n4430), .Z(n4437) );
  COND3X1 U3536 ( .A(n4438), .B(n4437), .C(n4436), .D(n4435), .Z(n853) );
  CIVX2 U3537 ( .A(n4441), .Z(n4448) );
  COND3X1 U3538 ( .A(n4454), .B(n3208), .C(n4453), .D(n4452), .Z(n854) );
  CND2X1 U3539 ( .A(n4456), .B(n4455), .Z(n4465) );
  CND2IX1 U3540 ( .B(n4553), .A(n4461), .Z(n4464) );
  CND2IX1 U3541 ( .B(n4553), .A(n4468), .Z(n4473) );
  COND3X1 U3542 ( .A(n3409), .B(res_not_wire[42]), .C(n3211), .D(n4469), .Z(
        n4472) );
  CND2IX1 U3543 ( .B(n4486), .A(n4485), .Z(n842) );
  CIVX2 U3544 ( .A(n4488), .Z(n4489) );
  CENX1 U3545 ( .A(n114), .B(n4506), .Z(n4507) );
  CND2IX1 U3546 ( .B(n3496), .A(n4507), .Z(n4510) );
  CIVX2 U3547 ( .A(i[31]), .Z(n4513) );
  CMXI2X1 U3548 ( .A0(n4522), .A1(n4521), .S(n4520), .Z(n4523) );
  CND2IX1 U3549 ( .B(n4553), .A(n4523), .Z(n4526) );
  CMXI2X1 U3550 ( .A0(n3508), .A1(n3505), .S(result[34]), .Z(n4528) );
  CEOX2 U3551 ( .A(n4533), .B(n4532), .Z(n4541) );
  CANR4CX1 U3552 ( .A(n4537), .B(res_not_wire[54]), .C(n4536), .D(n4535), .Z(
        n4540) );
  CND2IX1 U3553 ( .B(n4538), .A(n3200), .Z(n4539) );
  CND2IX1 U3554 ( .B(n4543), .A(n4542), .Z(n874) );
  CENX1 U3555 ( .A(n116), .B(n4548), .Z(n4549) );
  CND2IX1 U3556 ( .B(n3496), .A(n4549), .Z(n4552) );
  CMXI2X1 U3557 ( .A0(n3508), .A1(n3505), .S(result[55]), .Z(n4555) );
  CND2IX1 U3558 ( .B(n4556), .A(n2565), .Z(n891) );
  CND2IX1 U3559 ( .B(n4557), .A(n2562), .Z(n894) );
  CND2IX1 U3560 ( .B(n4558), .A(n2561), .Z(n895) );
  CND2IX1 U3561 ( .B(n4559), .A(n2555), .Z(n901) );
  CND2IX1 U3562 ( .B(n4560), .A(n2552), .Z(n904) );
  CIVX2 U3563 ( .A(n4564), .Z(n4563) );
  CMXI2X1 U3564 ( .A0(i[7]), .A1(n4565), .S(i[6]), .Z(n4568) );
  CIVX2 U3565 ( .A(n4579), .Z(n4577) );
  CND2IX1 U3566 ( .B(n4588), .A(n4587), .Z(n4592) );
  CND2IX1 U3567 ( .B(i[12]), .A(n4649), .Z(n4590) );
  CMXI2X1 U3568 ( .A0(i[15]), .A1(n4595), .S(i[14]), .Z(n4598) );
  CIVX2 U3569 ( .A(n4603), .Z(n4600) );
  CIVX2 U3570 ( .A(n4601), .Z(n4602) );
  CMXI2X1 U3571 ( .A0(n4605), .A1(n4604), .S(n3266), .Z(n935) );
  CND2IX1 U3572 ( .B(i[20]), .A(n4649), .Z(n4612) );
  CIVX2 U3573 ( .A(n4616), .Z(n4615) );
  CMXI2X1 U3574 ( .A0(i[23]), .A1(n4617), .S(i[22]), .Z(n4620) );
  CND2IX1 U3575 ( .B(i[24]), .A(n4649), .Z(n4628) );
  CIVX2 U3576 ( .A(n4640), .Z(n4633) );
  CMXI2X1 U3577 ( .A0(n4636), .A1(n2284), .S(i[27]), .Z(n4639) );
endmodule


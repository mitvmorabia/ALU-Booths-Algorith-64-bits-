
module multiplier ( result, valid, opera1, opera2, muordi, clock, reset, start
 );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input muordi, clock, reset, start;
  output valid;
  wire   opera2_63, N34, n52, n53, n55, n56, n100, n108, n110, n112, n114,
         n116, n118, n122, n124, n126, n128, n130, n132, n134, n136, n138,
         n140, n142, n144, n146, n148, n150, n152, n154, n156, n158, n160,
         n162, n164, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n1026, n1048, n1073, n1081, n1106, n1982, n1983, n1984,
         n1986, n1987, n1989, n1990, n1997, n1998, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2013, n2018,
         n2020, n2024, n2035, n2046, n2047, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2083, n2086, n2087, n2088, n2089,
         n2091, n2092, n2093, n2094, n2095, n2096, n2099, n2101, n2102, n2106,
         n2116, n2118, n2120, n2123, n2125, n2128, n2131, n2135, n2136, n2137,
         n2138, n2144, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2157, n2158, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2250, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2285, n2286, n2288, n2292, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2640, n2641, n2642, n2645, n2646, n2648,
         n2650, n2651, n2652, n2655, n2657, n2658, n2659, n2662, n2664, n2665,
         n2667, n2669, n2670, n2671, n2674, n2676, n2677, n2678, n2681, n2683,
         n2684, n2686, n2688, n2689, n2690, n2693, n2695, n2696, n2697, n2700,
         n2702, n2703, n2705, n2707, n2708, n2709, n2712, n2714, n2715, n2716,
         n2719, n2721, n2722, n2724, n2726, n2727, n2728, n2731, n2733, n2734,
         n2735, n2738, n2740, n2741, n2743, n2745, n2746, n2747, n2750, n2752,
         n2753, n2754, n2757, n2759, n2760, n2762, n2764, n2765, n2766, n2769,
         n2771, n2772, n2773, n2776, n2778, n2779, n2781, n2783, n2784, n2785,
         n2788, n2790, n2791, n2792, n2795, n2797, n2798, n2800, n2802, n2803,
         n2804, n2807, n2809, n2810, n2811, n2814, n2816, n2817, n2819, n2821,
         n2822, n2823, n2826, n2828, n2829, n2830, n2833, n2835, n2840, n2841,
         n2842, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2881, n2882, n2883, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769;
  wire   [63:0] res_not_wire;
  wire   [2:0] nst;
  wire   [31:0] i;
  tri   c_inop1;
  tri   c_inop2;
  tri   c_inres;
  assign opera2_63 = opera2[63];

  CTSX2 A5 ( .A(1'b1), .E(n1048), .Z(c_inres) );
  CTSX2 A4 ( .A(1'b0), .E(n1983), .Z(c_inop2) );
  CTSX2 A3 ( .A(1'b1), .E(opera2_63), .Z(c_inop2) );
  CTSX2 A6 ( .A(1'b0), .E(n100), .Z(c_inres) );
  CND2X2 U1545 ( .A(n2754), .B(n2760), .Z(n2765) );
  CAN3X2 U1624 ( .A(i[14]), .B(n2008), .C(i[15]), .Z(n2215) );
  CIVX2 U1684 ( .A(n2202), .Z(n1986) );
  CIVX2 U1685 ( .A(n2213), .Z(n1987) );
  CIVX2 U1687 ( .A(n2170), .Z(n1989) );
  CIVX2 U1688 ( .A(n2166), .Z(n1990) );
  CIVX2 U1695 ( .A(reset), .Z(n1997) );
  CIVX2 U1696 ( .A(n2157), .Z(n1998) );
  CIVX2 U1700 ( .A(n2218), .Z(n2002) );
  CIVX2 U1701 ( .A(n2217), .Z(n2003) );
  CIVX2 U1702 ( .A(n2243), .Z(n2004) );
  CIVX2 U1703 ( .A(n2209), .Z(n2005) );
  CIVX2 U1704 ( .A(i[18]), .Z(n2006) );
  CIVX2 U1705 ( .A(n2204), .Z(n2007) );
  CIVX2 U1706 ( .A(n2196), .Z(n2008) );
  CIVX2 U1707 ( .A(n2191), .Z(n2009) );
  CIVX2 U1709 ( .A(i[8]), .Z(n2011) );
  CIVX2 U1711 ( .A(res_not_wire[58]), .Z(n2013) );
  CIVX2 U1716 ( .A(res_not_wire[62]), .Z(n2018) );
  CIVX2 U1718 ( .A(n1081), .Z(n2020) );
  CIVX2 U1722 ( .A(n1073), .Z(n2024) );
  CIVX2 U1733 ( .A(result[41]), .Z(n2035) );
  CIVX2 U1744 ( .A(result[35]), .Z(n2046) );
  CIVX2 U1747 ( .A(result[29]), .Z(n2049) );
  CIVX2 U1748 ( .A(result[27]), .Z(n2050) );
  CIVX2 U1749 ( .A(result[25]), .Z(n2051) );
  CIVX2 U1750 ( .A(result[23]), .Z(n2052) );
  CIVX2 U1751 ( .A(result[21]), .Z(n2053) );
  CIVX2 U1752 ( .A(result[19]), .Z(n2054) );
  CIVX2 U1753 ( .A(result[17]), .Z(n2055) );
  CIVX2 U1754 ( .A(result[15]), .Z(n2056) );
  CIVX2 U1755 ( .A(result[13]), .Z(n2057) );
  CIVX2 U1756 ( .A(result[11]), .Z(n2058) );
  CIVX2 U1757 ( .A(result[9]), .Z(n2059) );
  CIVX2 U1758 ( .A(result[7]), .Z(n2060) );
  CIVX2 U1759 ( .A(result[5]), .Z(n2061) );
  CIVX2 U1760 ( .A(result[3]), .Z(n2062) );
  CIVX2 U1761 ( .A(result[1]), .Z(n2063) );
  CIVX2 U1762 ( .A(result[30]), .Z(n2064) );
  CIVX2 U1763 ( .A(result[28]), .Z(n2065) );
  CIVX2 U1764 ( .A(result[26]), .Z(n2066) );
  CIVX2 U1765 ( .A(result[24]), .Z(n2067) );
  CIVX2 U1766 ( .A(result[22]), .Z(n2068) );
  CIVX2 U1767 ( .A(result[20]), .Z(n2069) );
  CIVX2 U1768 ( .A(result[18]), .Z(n2070) );
  CIVX2 U1769 ( .A(result[16]), .Z(n2071) );
  CIVX2 U1770 ( .A(result[14]), .Z(n2072) );
  CIVX2 U1771 ( .A(result[12]), .Z(n2073) );
  CIVX2 U1772 ( .A(result[10]), .Z(n2074) );
  CIVX2 U1773 ( .A(result[8]), .Z(n2075) );
  CIVX2 U1774 ( .A(result[6]), .Z(n2076) );
  CIVX2 U1775 ( .A(result[4]), .Z(n2077) );
  CIVX2 U1776 ( .A(result[2]), .Z(n2078) );
  CIVX2 U1784 ( .A(n2181), .Z(n2086) );
  CIVX2 U1787 ( .A(i[0]), .Z(n2089) );
  CIVX2 U1789 ( .A(i[1]), .Z(n2091) );
  CIVX2 U1790 ( .A(i[24]), .Z(n2092) );
  CIVX2 U1791 ( .A(i[28]), .Z(n2093) );
  CIVX2 U1792 ( .A(i[29]), .Z(n2094) );
  CIVX2 U1793 ( .A(i[26]), .Z(n2095) );
  CIVX2 U1799 ( .A(n2842), .Z(n2101) );
  CIVX2 U1800 ( .A(n53), .Z(n2102) );
  CIVX2 U1816 ( .A(res_not_wire[4]), .Z(n2118) );
  CIVX2 U1821 ( .A(res_not_wire[8]), .Z(n2123) );
  CIVX2 U1823 ( .A(res_not_wire[52]), .Z(n2125) );
  CIVX2 U1826 ( .A(res_not_wire[46]), .Z(n2128) );
  CIVX2 U1829 ( .A(res_not_wire[28]), .Z(n2131) );
  CIVX2 U1844 ( .A(result[31]), .Z(n2146) );
  CIVX2 U1845 ( .A(i[21]), .Z(n2147) );
  CIVX2 U1847 ( .A(i[16]), .Z(n2149) );
  CIVX2 U1848 ( .A(i[14]), .Z(n2150) );
  CIVX2 U1849 ( .A(i[12]), .Z(n2151) );
  CIVX2 U1850 ( .A(i[10]), .Z(n2152) );
  CIVX2 U1851 ( .A(i[6]), .Z(n2153) );
  CAOR2X1 U1853 ( .A(i[31]), .B(n1989), .C(n2902), .D(n3059), .Z(n955) );
  COR4X1 U1856 ( .A(n2011), .B(n3060), .C(i[9]), .D(n2181), .Z(n2185) );
  COR4X1 U1858 ( .A(n2151), .B(n3060), .C(i[13]), .D(n2191), .Z(n2195) );
  COR4X1 U1860 ( .A(n3060), .B(n2204), .C(i[19]), .D(n2006), .Z(n2208) );
  CND2IX1 U1861 ( .B(n2211), .A(i[20]), .Z(n2210) );
  COR4X1 U1863 ( .A(n2095), .B(n3060), .C(i[27]), .D(n2223), .Z(n2227) );
  CAOR2X1 U1864 ( .A(valid), .B(n2885), .C(n3058), .D(n3768), .Z(n923) );
  CAN4X1 U1865 ( .A(n2238), .B(n2240), .C(n2241), .D(n2242), .Z(n2157) );
  CAN4X1 U1893 ( .A(i[21]), .B(i[20]), .C(i[22]), .D(n2847), .Z(n2217) );
  CAN4X1 U1894 ( .A(i[19]), .B(i[18]), .C(i[17]), .D(i[16]), .Z(n2847) );
  CAN4X1 U1895 ( .A(n56), .B(n53), .C(n1106), .D(reset), .Z(n2244) );
  CNR8X1 U1896 ( .A(i[1]), .B(i[19]), .C(i[16]), .D(i[2]), .E(n2849), .F(n2850), .G(n2846), .H(n2851), .Z(n2243) );
  COR6X1 U1898 ( .A(i[11]), .B(n2852), .C(n2850), .D(i[5]), .E(i[19]), .F(
        i[16]), .Z(n2853) );
  COR8X1 U1899 ( .A(i[20]), .B(i[17]), .C(i[22]), .D(i[21]), .E(i[26]), .F(
        i[24]), .G(i[9]), .H(i[30]), .Z(n2852) );
  COR8X1 U1900 ( .A(i[13]), .B(i[12]), .C(i[10]), .D(n2854), .E(i[28]), .F(
        i[27]), .G(i[25]), .H(n2855), .Z(n2850) );
  COR4X1 U1901 ( .A(i[29]), .B(i[6]), .C(i[7]), .D(i[8]), .Z(n2855) );
  COR4X1 U1902 ( .A(i[14]), .B(i[15]), .C(i[18]), .D(i[23]), .Z(n2854) );
  CND2IX1 U1903 ( .B(n2927), .A(nst[1]), .Z(n52) );
  CFD1X1 \res_not_reg[7]  ( .D(n912), .CP(clock), .Q(n3039), .QN(n158) );
  CFD1X1 \res_not_reg[9]  ( .D(n910), .CP(clock), .Q(n3037), .QN(n156) );
  CFD1QXL \res_not_reg[4]  ( .D(n915), .CP(clock), .Q(res_not_wire[4]) );
  CFD1QXL \nst_reg[2]  ( .D(n921), .CP(clock), .Q(nst[2]) );
  CFD1XL \res_not_reg[60]  ( .D(n859), .CP(clock), .Q(res_not_wire[60]), .QN(
        n3015) );
  CFD1QXL \nst_reg[0]  ( .D(n2909), .CP(clock), .Q(nst[0]) );
  CFD1QXL \result_reg[19]  ( .D(n806), .CP(clock), .Q(result[19]) );
  CFD1QXL \result_reg[1]  ( .D(n824), .CP(clock), .Q(result[1]) );
  CFD1QXL \result_reg[3]  ( .D(n822), .CP(clock), .Q(result[3]) );
  CFD1QXL \result_reg[2]  ( .D(n2911), .CP(clock), .Q(result[2]) );
  CFD1QXL \result_reg[29]  ( .D(n796), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[27]  ( .D(n798), .CP(clock), .Q(result[27]) );
  CFD1QXL \result_reg[25]  ( .D(n800), .CP(clock), .Q(result[25]) );
  CFD1QXL \result_reg[23]  ( .D(n802), .CP(clock), .Q(result[23]) );
  CFD1QXL \result_reg[21]  ( .D(n804), .CP(clock), .Q(result[21]) );
  CFD1QXL \result_reg[17]  ( .D(n808), .CP(clock), .Q(result[17]) );
  CFD1QXL \result_reg[15]  ( .D(n810), .CP(clock), .Q(result[15]) );
  CFD1QXL \result_reg[13]  ( .D(n812), .CP(clock), .Q(result[13]) );
  CFD1QXL \result_reg[11]  ( .D(n814), .CP(clock), .Q(result[11]) );
  CFD1QXL \result_reg[9]  ( .D(n816), .CP(clock), .Q(result[9]) );
  CFD1QXL \result_reg[7]  ( .D(n818), .CP(clock), .Q(result[7]) );
  CFD1QXL \result_reg[5]  ( .D(n820), .CP(clock), .Q(result[5]) );
  CFD1QXL \result_reg[30]  ( .D(n795), .CP(clock), .Q(result[30]) );
  CFD1QXL \result_reg[28]  ( .D(n797), .CP(clock), .Q(result[28]) );
  CFD1QXL \result_reg[26]  ( .D(n2913), .CP(clock), .Q(result[26]) );
  CFD1QXL \result_reg[24]  ( .D(n801), .CP(clock), .Q(result[24]) );
  CFD1QXL \result_reg[22]  ( .D(n803), .CP(clock), .Q(result[22]) );
  CFD1QXL \result_reg[20]  ( .D(n805), .CP(clock), .Q(result[20]) );
  CFD1QXL \result_reg[18]  ( .D(n807), .CP(clock), .Q(result[18]) );
  CFD1QXL \result_reg[16]  ( .D(n809), .CP(clock), .Q(result[16]) );
  CFD1QXL \result_reg[14]  ( .D(n811), .CP(clock), .Q(result[14]) );
  CFD1QXL \result_reg[12]  ( .D(n813), .CP(clock), .Q(result[12]) );
  CFD1QXL \result_reg[10]  ( .D(n815), .CP(clock), .Q(result[10]) );
  CFD1QXL \result_reg[8]  ( .D(n817), .CP(clock), .Q(result[8]) );
  CFD1QXL \result_reg[6]  ( .D(n819), .CP(clock), .Q(result[6]) );
  CFD1QXL \result_reg[4]  ( .D(n821), .CP(clock), .Q(result[4]) );
  CFD1QXL \result_reg[63]  ( .D(n919), .CP(clock), .Q(result[63]) );
  CFD1QXL \result_reg[0]  ( .D(n825), .CP(clock), .Q(result[0]) );
  CFD1QXL \res_not_reg[54]  ( .D(n865), .CP(clock), .Q(res_not_wire[54]) );
  CFD1QXL \res_not_reg[52]  ( .D(n867), .CP(clock), .Q(res_not_wire[52]) );
  CFD1XL \res_not_reg[53]  ( .D(n866), .CP(clock), .QN(n112) );
  CFD1XL \res_not_reg[57]  ( .D(n862), .CP(clock), .Q(n2955), .QN(n108) );
  CFD1XL \res_not_reg[55]  ( .D(n864), .CP(clock), .Q(n2903), .QN(n110) );
  CFD1XL \res_not_reg[51]  ( .D(n868), .CP(clock), .Q(n2861), .QN(n114) );
  CFD1XL \result_reg[59]  ( .D(n829), .CP(clock), .Q(result[59]), .QN(n3009)
         );
  CFD1XL \result_reg[61]  ( .D(n827), .CP(clock), .Q(result[61]), .QN(n2942)
         );
  CFD1QXL \res_not_reg[42]  ( .D(n877), .CP(clock), .Q(res_not_wire[42]) );
  CFD1XL \res_not_reg[45]  ( .D(n874), .CP(clock), .Q(n3697), .QN(n2872) );
  CFD1QXL \res_not_reg[48]  ( .D(n871), .CP(clock), .Q(res_not_wire[48]) );
  CFD1XL \res_not_reg[47]  ( .D(n872), .CP(clock), .Q(n2870), .QN(n118) );
  CFD1QXL \res_not_reg[50]  ( .D(n869), .CP(clock), .Q(res_not_wire[50]) );
  CFD1QXL \res_not_reg[46]  ( .D(n873), .CP(clock), .Q(res_not_wire[46]) );
  CFD1XL \res_not_reg[49]  ( .D(n870), .CP(clock), .Q(n2904), .QN(n116) );
  CFD1XL \result_reg[53]  ( .D(n835), .CP(clock), .Q(result[53]), .QN(n3003)
         );
  CFD1XL \result_reg[46]  ( .D(n842), .CP(clock), .Q(result[46]), .QN(n3026)
         );
  CFD1QXL \result_reg[45]  ( .D(n843), .CP(clock), .Q(result[45]) );
  CFD1XL \result_reg[55]  ( .D(n833), .CP(clock), .Q(result[55]), .QN(n3004)
         );
  CFD1XL \result_reg[57]  ( .D(n831), .CP(clock), .Q(result[57]), .QN(n3000)
         );
  CFD1QXL \result_reg[56]  ( .D(n832), .CP(clock), .Q(result[56]) );
  CFD1QXL \result_reg[54]  ( .D(n834), .CP(clock), .Q(result[54]) );
  CFD1QXL \result_reg[49]  ( .D(n839), .CP(clock), .Q(result[49]) );
  CFD1QXL \result_reg[48]  ( .D(n840), .CP(clock), .Q(result[48]) );
  CFD1QXL \res_not_reg[40]  ( .D(n879), .CP(clock), .Q(res_not_wire[40]) );
  CFD1XL \res_not_reg[43]  ( .D(n876), .CP(clock), .Q(n2901), .QN(n122) );
  CFD1QXL \i_reg[11]  ( .D(n943), .CP(clock), .Q(i[11]) );
  CFD1QXL \i_reg[31]  ( .D(n955), .CP(clock), .Q(i[31]) );
  CFD1XL \res_not_reg[39]  ( .D(n880), .CP(clock), .Q(n2937), .QN(n126) );
  CFD1XL \res_not_reg[41]  ( .D(n878), .CP(clock), .Q(n2869), .QN(n124) );
  CFD1XL \res_not_reg[37]  ( .D(n882), .CP(clock), .QN(n128) );
  CFD1QXL \res_not_reg[38]  ( .D(n881), .CP(clock), .Q(res_not_wire[38]) );
  CFD1QXL \i_reg[19]  ( .D(n935), .CP(clock), .Q(i[19]) );
  CFD1QXL \i_reg[16]  ( .D(n938), .CP(clock), .Q(i[16]) );
  CFD1QXL \result_reg[40]  ( .D(n848), .CP(clock), .Q(result[40]) );
  CFD1XL \result_reg[39]  ( .D(n849), .CP(clock), .Q(result[39]), .QN(n3018)
         );
  CFD1QXL \result_reg[43]  ( .D(n845), .CP(clock), .Q(result[43]) );
  CFD1XL \result_reg[38]  ( .D(n850), .CP(clock), .Q(result[38]), .QN(n3006)
         );
  CFD1QXL \result_reg[36]  ( .D(n852), .CP(clock), .Q(result[36]) );
  CFD1XL \result_reg[37]  ( .D(n851), .CP(clock), .Q(result[37]), .QN(n3002)
         );
  CFD1QXL \result_reg[42]  ( .D(n846), .CP(clock), .Q(result[42]) );
  CFD1XL \result_reg[51]  ( .D(n837), .CP(clock), .Q(result[51]), .QN(n3008)
         );
  CFD1XL \result_reg[50]  ( .D(n838), .CP(clock), .Q(result[50]), .QN(n3005)
         );
  CFD1QXL \result_reg[52]  ( .D(n836), .CP(clock), .Q(result[52]) );
  CFD1QXL \i_reg[30]  ( .D(n924), .CP(clock), .Q(i[30]) );
  CFD1QXL \res_not_reg[6]  ( .D(n913), .CP(clock), .Q(res_not_wire[6]) );
  CFD1QXL \i_reg[22]  ( .D(n932), .CP(clock), .Q(i[22]) );
  CFD1QXL \i_reg[25]  ( .D(n929), .CP(clock), .Q(i[25]) );
  CFD1QXL \i_reg[13]  ( .D(n941), .CP(clock), .Q(i[13]) );
  CFD1QXL \i_reg[17]  ( .D(n937), .CP(clock), .Q(i[17]) );
  CFD1QXL \i_reg[28]  ( .D(n926), .CP(clock), .Q(i[28]) );
  CFD1QXL \i_reg[29]  ( .D(n925), .CP(clock), .Q(i[29]) );
  CFD1XL \res_not_reg[15]  ( .D(n2915), .CP(clock), .Q(n3522), .QN(n150) );
  CFD1XL \res_not_reg[33]  ( .D(n886), .CP(clock), .Q(n3748), .QN(n132) );
  CFD1XL \res_not_reg[5]  ( .D(n914), .CP(clock), .Q(n2967), .QN(n160) );
  CFD1QXL \i_reg[23]  ( .D(n931), .CP(clock), .Q(i[23]) );
  CFD1XL \res_not_reg[35]  ( .D(n884), .CP(clock), .QN(n130) );
  CFD1QXL \res_not_reg[26]  ( .D(n893), .CP(clock), .Q(res_not_wire[26]) );
  CFD1QXL \res_not_reg[34]  ( .D(n885), .CP(clock), .Q(res_not_wire[34]) );
  CFD1XL \res_not_reg[13]  ( .D(n2916), .CP(clock), .Q(n3516), .QN(n152) );
  CFD1XL \res_not_reg[25]  ( .D(n2917), .CP(clock), .Q(n3553), .QN(n140) );
  CFD1XL \res_not_reg[27]  ( .D(n892), .CP(clock), .Q(n2966), .QN(n138) );
  CFD1QXL \i_reg[10]  ( .D(n944), .CP(clock), .Q(i[10]) );
  CFD1QXL \i_reg[6]  ( .D(n948), .CP(clock), .Q(i[6]) );
  CFD1QXL \i_reg[24]  ( .D(n930), .CP(clock), .Q(i[24]) );
  CFD1QXL \result_reg[32]  ( .D(n856), .CP(clock), .Q(result[32]) );
  CFD1XL \res_not_reg[31]  ( .D(n888), .CP(clock), .QN(n134) );
  CFD1QXL \res_not_reg[16]  ( .D(n903), .CP(clock), .Q(res_not_wire[16]) );
  CFD1XL \res_not_reg[23]  ( .D(n896), .CP(clock), .Q(n2965), .QN(n142) );
  CFD1QXL \i_reg[7]  ( .D(n947), .CP(clock), .Q(i[7]) );
  CFD1QXL \i_reg[9]  ( .D(n945), .CP(clock), .Q(i[9]) );
  CFD1QXL \i_reg[8]  ( .D(n946), .CP(clock), .Q(i[8]) );
  CFD1QXL \i_reg[12]  ( .D(n942), .CP(clock), .Q(i[12]) );
  CFD1QXL \i_reg[20]  ( .D(n934), .CP(clock), .Q(i[20]) );
  CFD1QXL \i_reg[27]  ( .D(n927), .CP(clock), .Q(i[27]) );
  CFD1QXL \i_reg[26]  ( .D(n928), .CP(clock), .Q(i[26]) );
  CTSX2 A1 ( .A(1'b1), .E(opera1[31]), .Z(c_inop1) );
  CTSX2 A2 ( .A(1'b0), .E(n2950), .Z(c_inop1) );
  CFD1XL \res_not_reg[17]  ( .D(n902), .CP(clock), .Q(n2905), .QN(n148) );
  CFD1XL \res_not_reg[22]  ( .D(n897), .CP(clock), .Q(res_not_wire[22]), .QN(
        n3028) );
  CFD1QXL \i_reg[15]  ( .D(n939), .CP(clock), .Q(i[15]) );
  CFD1QXL \i_reg[18]  ( .D(n936), .CP(clock), .Q(i[18]) );
  CFD1QX1 \res_not_reg[0]  ( .D(n2919), .CP(clock), .Q(res_not_wire[0]) );
  CFD1QXL \i_reg[3]  ( .D(n954), .CP(clock), .Q(i[3]) );
  CFD1QXL \res_not_reg[12]  ( .D(n907), .CP(clock), .Q(res_not_wire[12]) );
  CFD1XL \res_not_reg[24]  ( .D(n895), .CP(clock), .Q(res_not_wire[24]), .QN(
        n3027) );
  CFD1QXL \res_not_reg[18]  ( .D(n901), .CP(clock), .Q(res_not_wire[18]) );
  CFD1QXL \i_reg[4]  ( .D(n949), .CP(clock), .Q(i[4]) );
  CFD1XL \res_not_reg[3]  ( .D(n916), .CP(clock), .Q(n2862), .QN(n162) );
  CFD1QXL \i_reg[5]  ( .D(n953), .CP(clock), .Q(i[5]) );
  CFD1QXL \result_reg[31]  ( .D(n794), .CP(clock), .Q(result[31]) );
  CFD1QXL \i_reg[2]  ( .D(n950), .CP(clock), .Q(i[2]) );
  CFD1QXL \i_reg[1]  ( .D(n951), .CP(clock), .Q(i[1]) );
  CFD1QX1 \res_not_reg[30]  ( .D(n2924), .CP(clock), .Q(res_not_wire[30]) );
  CFD1QX1 \res_not_reg[28]  ( .D(n2925), .CP(clock), .Q(res_not_wire[28]) );
  CFD1QXL \result_reg[58]  ( .D(n830), .CP(clock), .Q(result[58]) );
  CFD4QXL \cst_reg[0]  ( .D(n55), .CP(clock), .SD(n1997), .Q(n56) );
  CFD4QXL \cst_reg[1]  ( .D(n52), .CP(clock), .SD(n1997), .Q(n53) );
  CFD2XL \cst_reg[2]  ( .D(N34), .CP(clock), .CD(n1997), .Q(n3764), .QN(n1106)
         );
  CFD1X1 \res_not_reg[29]  ( .D(n2928), .CP(clock), .Q(n3565), .QN(n136) );
  CFD1QXL valid_reg ( .D(n923), .CP(clock), .Q(valid) );
  CFD1QXL \i_reg[21]  ( .D(n933), .CP(clock), .Q(i[21]) );
  CFD1QXL \res_not_reg[32]  ( .D(n887), .CP(clock), .Q(res_not_wire[32]) );
  CFD1QXL \res_not_reg[44]  ( .D(n875), .CP(clock), .Q(res_not_wire[44]) );
  CFD1QXL \res_not_reg[56]  ( .D(n863), .CP(clock), .Q(res_not_wire[56]) );
  CFD1QXL \res_not_reg[36]  ( .D(n883), .CP(clock), .Q(res_not_wire[36]) );
  CFD1QXL \res_not_reg[63]  ( .D(n793), .CP(clock), .Q(n1026) );
  CFD1QXL \res_not_reg[62]  ( .D(n857), .CP(clock), .Q(res_not_wire[62]) );
  CFD1QXL \res_not_reg[61]  ( .D(n858), .CP(clock), .Q(n1081) );
  CFD1QXL \res_not_reg[59]  ( .D(n860), .CP(clock), .Q(n1073) );
  CFD1QXL \res_not_reg[58]  ( .D(n861), .CP(clock), .Q(res_not_wire[58]) );
  CFD1QXL \result_reg[33]  ( .D(n855), .CP(clock), .Q(result[33]) );
  CFD1QXL \result_reg[60]  ( .D(n828), .CP(clock), .Q(result[60]) );
  CFD1QXL \result_reg[44]  ( .D(n844), .CP(clock), .Q(result[44]) );
  CFD1QXL \result_reg[34]  ( .D(n854), .CP(clock), .Q(result[34]) );
  CFD1QXL \result_reg[47]  ( .D(n841), .CP(clock), .Q(result[47]) );
  CFD1QXL \result_reg[41]  ( .D(n847), .CP(clock), .Q(result[41]) );
  CFD1QXL \result_reg[35]  ( .D(n853), .CP(clock), .Q(result[35]) );
  CFD1XL \nst_reg[1]  ( .D(n2930), .CP(clock), .Q(nst[1]), .QN(n2047) );
  CFD1X1 sign_reg ( .D(n2931), .CP(clock), .Q(n1048), .QN(n100) );
  CFD1QXL \res_not_reg[2]  ( .D(n917), .CP(clock), .Q(res_not_wire[2]) );
  CFD1QXL \res_not_reg[14]  ( .D(n905), .CP(clock), .Q(res_not_wire[14]) );
  CFD1XL \res_not_reg[11]  ( .D(n2918), .CP(clock), .Q(n2895), .QN(n154) );
  CFD1XL \res_not_reg[1]  ( .D(n918), .CP(clock), .QN(n164) );
  CFD1QX1 \res_not_reg[8]  ( .D(n2922), .CP(clock), .Q(res_not_wire[8]) );
  CFD1X1 \res_not_reg[19]  ( .D(n2923), .CP(clock), .Q(n2876), .QN(n146) );
  CFD1QX1 \result_reg[62]  ( .D(n826), .CP(clock), .Q(result[62]) );
  CFD1QXL \i_reg[14]  ( .D(n940), .CP(clock), .Q(i[14]) );
  CFD1QX1 \res_not_reg[20]  ( .D(n2926), .CP(clock), .Q(res_not_wire[20]) );
  CFD1X1 \res_not_reg[21]  ( .D(n2856), .CP(clock), .QN(n144) );
  CFD1QXL \i_reg[0]  ( .D(n952), .CP(clock), .Q(i[0]) );
  CFD1QXL \res_not_reg[10]  ( .D(n909), .CP(clock), .Q(res_not_wire[10]) );
  COND3XL U1904 ( .A(n2640), .B(n2882), .C(n2641), .D(n2642), .Z(n825) );
  CNIVX1 U1905 ( .A(n898), .Z(n2856) );
  CND2X2 U1906 ( .A(n2735), .B(n2741), .Z(n2746) );
  COND1X1 U1907 ( .A(n3237), .B(n3247), .C(n3236), .Z(n3238) );
  CIVX1 U1908 ( .A(n3164), .Z(n3128) );
  CND2XL U1909 ( .A(result[43]), .B(n3128), .Z(n3165) );
  CNR3X4 U1910 ( .A(n2772), .B(n2766), .C(n2765), .Z(n2773) );
  CANR1X1 U1911 ( .A(n3365), .B(n3155), .C(result[34]), .Z(n3156) );
  CEOX2 U1912 ( .A(opera1[7]), .B(opera1[31]), .Z(n2992) );
  CND2XL U1913 ( .A(result[44]), .B(n2969), .Z(n3169) );
  CND2X1 U1914 ( .A(n3110), .B(n3109), .Z(n3233) );
  CENXL U1915 ( .A(n2888), .B(n3667), .Z(n3669) );
  CND2X1 U1916 ( .A(n3160), .B(n3143), .Z(n3159) );
  CND2IX2 U1917 ( .B(n3113), .A(n3114), .Z(n3118) );
  CIVX1 U1918 ( .A(n2865), .Z(n3209) );
  COND2X2 U1919 ( .A(n3158), .B(n3159), .C(n3575), .D(n3574), .Z(n3264) );
  CANR5CX2 U1920 ( .A(result[35]), .B(n2970), .C(n3585), .Z(n3575) );
  CNR4X2 U1921 ( .A(n3099), .B(n3117), .C(n3176), .D(n3153), .Z(n3100) );
  CND3X2 U1922 ( .A(n2951), .B(n3098), .C(c_inop1), .Z(n3153) );
  CND2IX1 U1923 ( .B(n3239), .A(n3238), .Z(n3241) );
  CND2X1 U1924 ( .A(n3653), .B(n3654), .Z(n3665) );
  CNR2X1 U1925 ( .A(n3088), .B(n148), .Z(n3042) );
  COND4CX1 U1926 ( .A(n3171), .B(n3279), .C(n3170), .D(n3169), .Z(n3645) );
  COND1XL U1927 ( .A(n3287), .B(n3285), .C(n2995), .Z(n3170) );
  CND2XL U1928 ( .A(n3289), .B(n3013), .Z(n3648) );
  CND2X1 U1929 ( .A(n3381), .B(n3380), .Z(n3702) );
  CND2IX1 U1930 ( .B(n3240), .A(n3241), .Z(n3381) );
  CENX1 U1931 ( .A(n3610), .B(n3611), .Z(n3614) );
  CEOX1 U1932 ( .A(n3714), .B(n3713), .Z(n2962) );
  CENX1 U1933 ( .A(n3702), .B(n3701), .Z(n3703) );
  CND2X1 U1934 ( .A(res_not_wire[6]), .B(n3074), .Z(n3426) );
  CIVX2 U1935 ( .A(opera1[31]), .Z(n2950) );
  CIVX3 U1936 ( .A(opera2_63), .Z(n1983) );
  COR3X1 U1937 ( .A(n3107), .B(n3103), .C(n3378), .Z(n3386) );
  CND2IX1 U1938 ( .B(n3610), .A(n3611), .Z(n3620) );
  CIVXL U1939 ( .A(n2863), .Z(n3611) );
  CANR1XL U1940 ( .A(n3166), .B(n3111), .C(n2857), .Z(n2969) );
  CIVX2 U1941 ( .A(n3167), .Z(n2857) );
  CND2IX1 U1942 ( .B(n3319), .A(n2944), .Z(n3225) );
  COR2XL U1943 ( .A(n3426), .B(n3075), .Z(n3510) );
  CNR2X1 U1944 ( .A(n3158), .B(n3047), .Z(n3266) );
  CNR2X1 U1945 ( .A(n3121), .B(n3153), .Z(n2971) );
  COND1XL U1946 ( .A(n3177), .B(n3102), .C(n3214), .Z(n3207) );
  CEOX1 U1947 ( .A(n2993), .B(n3160), .Z(n3161) );
  CND2IX1 U1948 ( .B(n3133), .A(result[42]), .Z(n3278) );
  CND2IX1 U1949 ( .B(n3681), .A(res_not_wire[54]), .Z(n3336) );
  CAOR1XL U1950 ( .A(n3039), .B(n3500), .C(res_not_wire[8]), .Z(n3430) );
  CNR2X1 U1951 ( .A(n3006), .B(n3046), .Z(n3735) );
  CND2IX1 U1952 ( .B(n3136), .A(result[40]), .Z(n3270) );
  CAN3X1 U1953 ( .A(n3218), .B(n2858), .C(n3339), .Z(n2896) );
  CIVX2 U1954 ( .A(n3346), .Z(n2858) );
  CENX1 U1955 ( .A(n3386), .B(n3385), .Z(n3396) );
  CND2IX1 U1956 ( .B(n3327), .A(n3205), .Z(n3323) );
  CND2IX1 U1957 ( .B(n3656), .A(n2890), .Z(n3658) );
  CND2X1 U1958 ( .A(n3691), .B(n3096), .Z(n3710) );
  CND4X1 U1959 ( .A(n2859), .B(res_not_wire[14]), .C(n3516), .D(n3522), .Z(
        n3088) );
  CIVX2 U1960 ( .A(n3076), .Z(n2859) );
  CEOXL U1961 ( .A(n122), .B(n3646), .Z(n3290) );
  CENX1 U1962 ( .A(n3199), .B(n3198), .Z(n3201) );
  CND2X1 U1963 ( .A(n3162), .B(n3163), .Z(n3279) );
  CND2X1 U1964 ( .A(n2862), .B(n3491), .Z(n3420) );
  CND2IX1 U1965 ( .B(n3206), .A(result[52]), .Z(n3326) );
  CND2X1 U1966 ( .A(n3093), .B(n2893), .Z(n3733) );
  CND3XL U1967 ( .A(n3679), .B(n2936), .C(res_not_wire[52]), .Z(n3681) );
  CENX1 U1968 ( .A(result[60]), .B(n3382), .Z(n2860) );
  CIVX2 U1969 ( .A(n2860), .Z(n3701) );
  CENXL U1970 ( .A(n2996), .B(n3712), .Z(n2973) );
  COR4X1 U1971 ( .A(n3426), .B(n3076), .C(n152), .D(n3036), .Z(n3523) );
  CNR2X1 U1972 ( .A(n2138), .B(n3046), .Z(n3307) );
  CND3XL U1973 ( .A(res_not_wire[28]), .B(res_not_wire[30]), .C(n3565), .Z(
        n3255) );
  CEOX1 U1974 ( .A(opera1[8]), .B(opera1[31]), .Z(n2991) );
  CND4X1 U1975 ( .A(n2937), .B(n3093), .C(n2893), .D(res_not_wire[40]), .Z(
        n3637) );
  COND1XL U1976 ( .A(n3148), .B(n3144), .C(n3149), .Z(n3738) );
  COND1XL U1977 ( .A(n3128), .B(result[43]), .C(n3165), .Z(n3280) );
  COND3X1 U1978 ( .A(n2863), .B(n3610), .C(n3621), .D(n3619), .Z(n3623) );
  COND1XL U1979 ( .A(n3340), .B(n3341), .C(n3339), .Z(n3345) );
  COND1XL U1980 ( .A(n3762), .B(n3404), .C(n3406), .Z(n3407) );
  CND2X1 U1981 ( .A(n2861), .B(n2934), .Z(n3328) );
  CND2IX1 U1982 ( .B(n3531), .A(res_not_wire[18]), .Z(n3454) );
  CND4X1 U1983 ( .A(n2862), .B(n3073), .C(n3491), .D(res_not_wire[4]), .Z(
        n3496) );
  COR2X1 U1984 ( .A(n3250), .B(n3249), .Z(n2864) );
  CMXI2X1 U1985 ( .A0(n3018), .A1(result[39]), .S(n3138), .Z(n3618) );
  CENX1 U1986 ( .A(n3110), .B(n3106), .Z(n3234) );
  CND4X1 U1987 ( .A(res_not_wire[46]), .B(n3697), .C(n3289), .D(n3013), .Z(
        n3601) );
  CAOR1X1 U1988 ( .A(n3153), .B(n3154), .C(result[33]), .Z(n3365) );
  CMXI2X1 U1989 ( .A0(n3009), .A1(result[59]), .S(n3105), .Z(n3240) );
  COR2X1 U1990 ( .A(n3637), .B(n124), .Z(n3639) );
  CANR2X1 U1991 ( .A(n3264), .B(n2866), .C(result[37]), .D(n2867), .Z(n2863)
         );
  CAN2X1 U1992 ( .A(n3342), .B(n3343), .Z(n3344) );
  CND2XL U1993 ( .A(n3015), .B(n3700), .Z(n3376) );
  CNR2X1 U1994 ( .A(n2942), .B(n3047), .Z(n3397) );
  CND2IX1 U1995 ( .B(n3567), .A(res_not_wire[30]), .Z(n3482) );
  CENX1 U1996 ( .A(n3039), .B(n3426), .Z(n3501) );
  COND3X1 U1997 ( .A(n2973), .B(n3044), .C(n2864), .D(n3252), .Z(n832) );
  CNR2IX1 U1998 ( .B(n3017), .A(n3119), .Z(n2985) );
  CNR3X1 U1999 ( .A(n3199), .B(n3198), .C(n3194), .Z(n2865) );
  CND2X1 U2000 ( .A(n3663), .B(n3204), .Z(n3202) );
  CND2IX1 U2001 ( .B(n3207), .A(result[48]), .Z(n3338) );
  COR2X1 U2002 ( .A(n134), .B(n3255), .Z(n3086) );
  CIVX2 U2003 ( .A(n3263), .Z(n2866) );
  CIVXL U2004 ( .A(n3161), .Z(n2867) );
  COR2X1 U2005 ( .A(n3601), .B(n118), .Z(n3603) );
  CND2IX1 U2006 ( .B(n3223), .A(result[49]), .Z(n3310) );
  CEOX1 U2007 ( .A(result[58]), .B(n3234), .Z(n3711) );
  CND2X1 U2008 ( .A(n2936), .B(res_not_wire[52]), .Z(n3678) );
  CIVDX1 U2009 ( .A(n3328), .Z0(n2936), .Z1(n2935) );
  CEOX1 U2010 ( .A(opera2[0]), .B(opera2_63), .Z(n2646) );
  CAOR1X1 U2011 ( .A(n3289), .B(n2901), .C(res_not_wire[44]), .Z(n3647) );
  CENX1 U2012 ( .A(result[40]), .B(n3136), .Z(n3011) );
  CND2IXL U2013 ( .B(n2941), .A(n3408), .Z(n2947) );
  CND4X1 U2014 ( .A(n2956), .B(n2955), .C(n1073), .D(res_not_wire[58]), .Z(
        n3700) );
  CND3XL U2015 ( .A(n3500), .B(n2905), .C(n3077), .Z(n3531) );
  CIVX2 U2016 ( .A(n3426), .Z(n3500) );
  CNR2X1 U2017 ( .A(n3004), .B(n3047), .Z(n3694) );
  CEOXL U2018 ( .A(n3302), .B(n3303), .Z(n3296) );
  CENX1 U2019 ( .A(n3209), .B(n3208), .Z(n3211) );
  COND4CXL U2020 ( .A(n2993), .B(n3140), .C(n3017), .D(n3141), .Z(n3142) );
  CMXI2X1 U2021 ( .A0(n3004), .A1(result[55]), .S(n3185), .Z(n3337) );
  CND2X1 U2022 ( .A(n3740), .B(result[32]), .Z(n3742) );
  CND2X1 U2023 ( .A(n3310), .B(n3673), .Z(n3321) );
  CENX1 U2024 ( .A(result[51]), .B(n3201), .Z(n2868) );
  CIVX2 U2025 ( .A(n2868), .Z(n3663) );
  CND3X1 U2026 ( .A(n2869), .B(res_not_wire[42]), .C(n3094), .Z(n3646) );
  CENX1 U2027 ( .A(opera2[2]), .B(opera2_63), .Z(n2658) );
  CANR5CXL U2028 ( .A(n3132), .B(result[41]), .C(n3634), .Z(n3635) );
  CEOXL U2029 ( .A(n3599), .B(n3341), .Z(n2975) );
  COR2X1 U2030 ( .A(n3747), .B(n132), .Z(n3750) );
  CND2IX1 U2031 ( .B(n3241), .A(n3240), .Z(n3242) );
  COR2X1 U2032 ( .A(n3733), .B(n126), .Z(n3043) );
  CND3X1 U2033 ( .A(n2870), .B(n3095), .C(res_not_wire[48]), .Z(n3656) );
  CND2IX1 U2034 ( .B(n3408), .A(n2941), .Z(n2948) );
  CNR2X1 U2035 ( .A(n3009), .B(n3048), .Z(n3705) );
  CAOR1X1 U2036 ( .A(n2876), .B(n3535), .C(res_not_wire[20]), .Z(n3455) );
  CND2X1 U2037 ( .A(n3027), .B(n3549), .Z(n3466) );
  COR4X1 U2038 ( .A(n3426), .B(n3075), .C(n154), .D(n2116), .Z(n3512) );
  COR2X1 U2039 ( .A(n3564), .B(n136), .Z(n3567) );
  CND2IX1 U2040 ( .B(n3178), .A(n3168), .Z(n3097) );
  COND1XL U2041 ( .A(n3126), .B(n2994), .C(n3166), .Z(n3164) );
  COND1XL U2042 ( .A(n3129), .B(n2992), .C(n3137), .Z(n3138) );
  CND2IX1 U2043 ( .B(n3222), .A(result[54]), .Z(n3343) );
  CMXI2X1 U2044 ( .A0(n3002), .A1(result[37]), .S(n3161), .Z(n3263) );
  CAN2X1 U2045 ( .A(n3225), .B(n3324), .Z(n3676) );
  CND4X1 U2046 ( .A(n2871), .B(res_not_wire[10]), .C(n2895), .D(
        res_not_wire[12]), .Z(n3076) );
  CIVX2 U2047 ( .A(n3075), .Z(n2871) );
  CND3XL U2048 ( .A(n3764), .B(n53), .C(n56), .Z(n3067) );
  CND2XL U2049 ( .A(n124), .B(n3637), .Z(n3638) );
  CND2XL U2050 ( .A(n118), .B(n3601), .Z(n3602) );
  CND2X1 U2051 ( .A(n132), .B(n3747), .Z(n3749) );
  CENX1 U2052 ( .A(n126), .B(n3733), .Z(n2998) );
  CENX1 U2053 ( .A(n3269), .B(n3634), .Z(n3273) );
  CND2X1 U2054 ( .A(n3310), .B(n3673), .Z(n3313) );
  CEOXL U2055 ( .A(n110), .B(n3336), .Z(n3692) );
  CANR2X2 U2056 ( .A(result[45]), .B(n3173), .C(n3172), .D(n3645), .Z(n3303)
         );
  CNR2X1 U2057 ( .A(n2872), .B(n3648), .Z(n3035) );
  CND2XL U2058 ( .A(n112), .B(n3678), .Z(n3680) );
  CNR2XL U2059 ( .A(n108), .B(n3710), .Z(n3016) );
  CAOR1X1 U2060 ( .A(res_not_wire[4]), .B(n3034), .C(n2967), .Z(n2907) );
  CEOX1 U2061 ( .A(n3541), .B(n144), .Z(n3542) );
  CND2IX1 U2062 ( .B(n3463), .A(n3465), .Z(n3549) );
  CND2X1 U2063 ( .A(n136), .B(n3564), .Z(n3566) );
  CMXI2X1 U2064 ( .A0(n100), .A1(n3591), .S(n2158), .Z(n956) );
  CAOR1X1 U2065 ( .A(n2947), .B(n2948), .C(n3044), .Z(n3399) );
  CIVDX1 U2066 ( .A(opera1[31]), .Z0(n2874), .Z1(n2873) );
  CEOXL U2067 ( .A(n3576), .B(n3575), .Z(n2974) );
  CND2X1 U2068 ( .A(res_not_wire[22]), .B(n3001), .Z(n3464) );
  CENX1 U2069 ( .A(n2963), .B(n2899), .Z(n3121) );
  CENX2 U2070 ( .A(opera1[1]), .B(opera1[31]), .Z(n3150) );
  CANR3X1 U2071 ( .A(n3592), .B(n2886), .C(n3190), .D(n3220), .Z(n3217) );
  CND2X1 U2072 ( .A(n3323), .B(n3326), .Z(n3319) );
  COND1X1 U2073 ( .A(n3600), .B(n3599), .C(n3338), .Z(n3311) );
  CND2IX1 U2074 ( .B(n2235), .A(n3752), .Z(n3066) );
  CANR1X1 U2075 ( .A(n3738), .B(n3157), .C(n3156), .Z(n3585) );
  CND3XL U2076 ( .A(result[34]), .B(n3365), .C(n3155), .Z(n3157) );
  CNR4X1 U2077 ( .A(n3464), .B(n3087), .C(n3086), .D(n3085), .Z(n3091) );
  CND3X1 U2078 ( .A(n3042), .B(n2964), .C(n3089), .Z(n3090) );
  CENX1 U2079 ( .A(n3593), .B(n3592), .Z(n3595) );
  CND2X1 U2080 ( .A(n3050), .B(n2683), .Z(n2681) );
  CAN3X2 U2081 ( .A(res_not_wire[20]), .B(n2876), .C(n3540), .Z(n2875) );
  CIVX2 U2082 ( .A(n3752), .Z(n3049) );
  CNIVX1 U2083 ( .A(n1983), .Z(n2877) );
  CND2XL U2084 ( .A(n3672), .B(n3671), .Z(n837) );
  CIVDX1 U2085 ( .A(opera1[31]), .Z0(n2879), .Z1(n2878) );
  CNR3X2 U2086 ( .A(n2696), .B(n2690), .C(n2689), .Z(n2697) );
  CND2X1 U2087 ( .A(n2678), .B(n2684), .Z(n2689) );
  CIVDX2 U2088 ( .A(n2250), .Z0(n2881), .Z1(n2882) );
  CND2IX1 U2089 ( .B(n3067), .A(n3752), .Z(n2250) );
  CIVX1 U2090 ( .A(n3066), .Z(n2883) );
  CEOX2 U2091 ( .A(opera1[31]), .B(opera1[0]), .Z(n2951) );
  COAN1X1 U2092 ( .A(n3147), .B(n3146), .C(n3145), .Z(n2970) );
  CENX1 U2093 ( .A(c_inop1), .B(n2951), .Z(n3069) );
  CAOR1X1 U2094 ( .A(n3065), .B(n3064), .C(n3063), .Z(n3752) );
  COND1X1 U2095 ( .A(n2233), .B(n3061), .C(i[31]), .Z(n3064) );
  CND2X1 U2096 ( .A(result[0]), .B(n2883), .Z(n3746) );
  CEOX1 U2097 ( .A(opera1[10]), .B(opera1[31]), .Z(n3012) );
  CENX1 U2098 ( .A(opera1[2]), .B(opera1[31]), .Z(n3120) );
  CIVX2 U2099 ( .A(opera1[3]), .Z(n2963) );
  CEOX1 U2100 ( .A(opera1[11]), .B(opera1[31]), .Z(n2994) );
  CEOX1 U2101 ( .A(opera1[6]), .B(opera1[31]), .Z(n3017) );
  CEOX1 U2102 ( .A(opera1[4]), .B(opera1[31]), .Z(n3010) );
  CEOX1 U2103 ( .A(opera1[5]), .B(opera1[31]), .Z(n2993) );
  CIVX2 U2104 ( .A(n3108), .Z(n2939) );
  CENX1 U2105 ( .A(opera1[12]), .B(opera1[31]), .Z(n3111) );
  CND2X1 U2106 ( .A(n2992), .B(n2991), .Z(n3113) );
  CND2X1 U2107 ( .A(n2994), .B(n3012), .Z(n3112) );
  CND2X1 U2108 ( .A(n2993), .B(n3010), .Z(n3119) );
  CIVX2 U2109 ( .A(n3111), .Z(n3168) );
  CIVX2 U2110 ( .A(n3208), .Z(n2940) );
  CIVX2 U2111 ( .A(n3120), .Z(n3148) );
  CIVX2 U2112 ( .A(n3150), .Z(n3098) );
  CEOX1 U2113 ( .A(result[56]), .B(n3229), .Z(n3220) );
  CNR2X1 U2114 ( .A(n2658), .B(n2651), .Z(n2968) );
  CND2X1 U2115 ( .A(c_inop2), .B(n2646), .Z(n2652) );
  CENX1 U2116 ( .A(n2942), .B(n3396), .Z(n3395) );
  CNR2X1 U2117 ( .A(n3235), .B(n3711), .Z(n3236) );
  CND2X1 U2118 ( .A(result[32]), .B(n3740), .Z(n3364) );
  CND3X1 U2119 ( .A(i[26]), .B(n2001), .C(i[27]), .Z(n2232) );
  CENX1 U2120 ( .A(n3142), .B(n3006), .Z(n3610) );
  COR2X1 U2121 ( .A(n3004), .B(n3185), .Z(n3686) );
  CIVX2 U2122 ( .A(n3336), .Z(n3691) );
  CENX1 U2123 ( .A(n3393), .B(n3405), .Z(n2941) );
  CND3X1 U2124 ( .A(n3037), .B(n3039), .C(res_not_wire[8]), .Z(n3075) );
  CND2X1 U2125 ( .A(n2716), .B(n2722), .Z(n2727) );
  CND2IX1 U2126 ( .B(n2803), .A(n2959), .Z(n2822) );
  CNR2X1 U2127 ( .A(n164), .B(n3415), .Z(n3072) );
  CND2X1 U2128 ( .A(res_not_wire[0]), .B(c_inres), .Z(n3486) );
  CNR2IX1 U2129 ( .B(n3740), .A(n3044), .Z(n3070) );
  CND2X1 U2130 ( .A(i[3]), .B(n2165), .Z(n2171) );
  CND3X1 U2131 ( .A(i[12]), .B(n2009), .C(i[13]), .Z(n2196) );
  CND3X1 U2132 ( .A(i[24]), .B(n2002), .C(i[25]), .Z(n2223) );
  CND3X1 U2133 ( .A(i[6]), .B(n2087), .C(i[7]), .Z(n2181) );
  CND3X1 U2134 ( .A(i[4]), .B(n2088), .C(i[5]), .Z(n2176) );
  CND3X1 U2135 ( .A(i[10]), .B(n2010), .C(i[11]), .Z(n2191) );
  CND3X1 U2136 ( .A(n2215), .B(n2217), .C(i[23]), .Z(n2218) );
  CIVX2 U2137 ( .A(n3646), .Z(n3289) );
  CND3X1 U2138 ( .A(i[8]), .B(n2086), .C(i[9]), .Z(n2186) );
  CAN2X1 U2139 ( .A(n2945), .B(n2946), .Z(n3713) );
  CND2X1 U2140 ( .A(n3402), .B(n3401), .Z(n3571) );
  CENX1 U2141 ( .A(res_not_wire[10]), .B(n3510), .Z(n3434) );
  CENX1 U2142 ( .A(n146), .B(n3535), .Z(n3536) );
  CENX1 U2143 ( .A(res_not_wire[0]), .B(c_inres), .Z(n2640) );
  CIVX2 U2144 ( .A(n3037), .Z(n3038) );
  COAN1X1 U2145 ( .A(n2235), .B(n2004), .C(n3062), .Z(n2885) );
  CIVDX1 U2146 ( .A(opera1[31]), .Z0(n2899), .Z1(n2900) );
  CAN2X1 U2147 ( .A(n3338), .B(n3304), .Z(n2886) );
  COR2X1 U2148 ( .A(n2101), .B(n3049), .Z(n2887) );
  CENX1 U2149 ( .A(result[52]), .B(n3206), .Z(n2888) );
  CNR2X1 U2150 ( .A(n2235), .B(n1989), .Z(n2161) );
  CNR2XL U2151 ( .A(n3117), .B(n3167), .Z(n2889) );
  CAN2X1 U2152 ( .A(res_not_wire[50]), .B(n2904), .Z(n2890) );
  CIVX2 U2153 ( .A(n3066), .Z(n2891) );
  CAN2X1 U2154 ( .A(n3082), .B(n3081), .Z(n2892) );
  CAN2X1 U2155 ( .A(res_not_wire[38]), .B(n3612), .Z(n2893) );
  CAN3X2 U2156 ( .A(n3343), .B(n3686), .C(n3342), .Z(n2894) );
  CAN3X2 U2157 ( .A(n2881), .B(n3747), .C(n3371), .Z(n2897) );
  CAN3X2 U2158 ( .A(n2881), .B(n3579), .C(n3578), .Z(n2898) );
  COAN1X1 U2159 ( .A(n2233), .B(n3061), .C(i[31]), .Z(n2902) );
  CNIVX1 U2160 ( .A(n2652), .Z(n2953) );
  COR2X1 U2161 ( .A(n2810), .B(n2804), .Z(n2906) );
  CNIVXL U2162 ( .A(muordi), .Z(n2933) );
  CNIVX1 U2163 ( .A(n3758), .Z(n2908) );
  CNIVX1 U2164 ( .A(n957), .Z(n2909) );
  CENXL U2165 ( .A(opera2[1]), .B(opera2_63), .Z(n2651) );
  CNIVX1 U2166 ( .A(n2664), .Z(n2910) );
  CNIVX1 U2167 ( .A(n823), .Z(n2911) );
  CND2X1 U2168 ( .A(n2828), .B(n3050), .Z(n2826) );
  CEOXL U2169 ( .A(opera2[27]), .B(opera2_63), .Z(n2817) );
  CENX1 U2170 ( .A(opera2[25]), .B(opera2_63), .Z(n2804) );
  CNIVX1 U2171 ( .A(n2804), .Z(n2912) );
  CEOXL U2172 ( .A(n2803), .B(n2912), .Z(n2802) );
  CND2X1 U2173 ( .A(n2676), .B(n3050), .Z(n2674) );
  CENXL U2174 ( .A(opera2[28]), .B(opera2_63), .Z(n2823) );
  CNIVX1 U2175 ( .A(n799), .Z(n2913) );
  CND2X1 U2176 ( .A(n3051), .B(n2797), .Z(n2795) );
  CEOXL U2177 ( .A(opera2[24]), .B(opera2_63), .Z(n2798) );
  CEOXL U2178 ( .A(opera2[21]), .B(opera2_63), .Z(n2779) );
  CENXL U2179 ( .A(opera2[22]), .B(opera2_63), .Z(n2785) );
  CENXL U2180 ( .A(opera2[19]), .B(opera2_63), .Z(n2766) );
  CND2X1 U2181 ( .A(n2771), .B(n3050), .Z(n2769) );
  CEOXL U2182 ( .A(opera2[18]), .B(opera2_63), .Z(n2760) );
  CEOXL U2183 ( .A(opera2[15]), .B(opera2_63), .Z(n2741) );
  CENXL U2184 ( .A(opera2[16]), .B(opera2_63), .Z(n2747) );
  CENXL U2185 ( .A(opera2[13]), .B(opera2_63), .Z(n2728) );
  CEOXL U2186 ( .A(opera2[12]), .B(opera2_63), .Z(n2722) );
  CEOXL U2187 ( .A(opera2[9]), .B(opera2_63), .Z(n2703) );
  CENXL U2188 ( .A(opera2[10]), .B(opera2_63), .Z(n2709) );
  CENXL U2189 ( .A(opera2[7]), .B(opera2_63), .Z(n2690) );
  CEOXL U2190 ( .A(opera2[6]), .B(opera2_63), .Z(n2684) );
  CENXL U2191 ( .A(opera2[4]), .B(opera2_63), .Z(n2671) );
  CNIVX1 U2192 ( .A(n2645), .Z(n2914) );
  CNIVX1 U2193 ( .A(n904), .Z(n2915) );
  CNIVX1 U2194 ( .A(n906), .Z(n2916) );
  CNIVX1 U2195 ( .A(n894), .Z(n2917) );
  COND1X1 U2196 ( .A(n142), .B(n3058), .C(n2274), .Z(n896) );
  CNIVX1 U2197 ( .A(n908), .Z(n2918) );
  CNIVX1 U2198 ( .A(n920), .Z(n2919) );
  CNIVXL U2199 ( .A(opera2[31]), .Z(n2921) );
  CND2X2 U2200 ( .A(n3083), .B(n2892), .Z(n794) );
  CIVDXL U2201 ( .A(opera2[30]), .Z0(n1984) );
  CNIVX1 U2202 ( .A(n911), .Z(n2922) );
  CIVXL U2203 ( .A(res_not_wire[10]), .Z(n2116) );
  CNIVX1 U2204 ( .A(n900), .Z(n2923) );
  CNIVX1 U2205 ( .A(n889), .Z(n2924) );
  CNIVX1 U2206 ( .A(n891), .Z(n2925) );
  CNIVX1 U2207 ( .A(n899), .Z(n2926) );
  CDLY1XL U2208 ( .A(start), .Z(n2927) );
  CNR2IXL U2209 ( .B(nst[2]), .A(n2927), .Z(N34) );
  CNIVX1 U2210 ( .A(n2929), .Z(n2928) );
  CNIVX1 U2211 ( .A(n890), .Z(n2929) );
  CNIVX1 U2212 ( .A(n922), .Z(n2930) );
  CNIVX1 U2213 ( .A(n2932), .Z(n2931) );
  CNIVX1 U2214 ( .A(n956), .Z(n2932) );
  CNR2XL U2215 ( .A(n2101), .B(n2933), .Z(n2158) );
  CIVX2 U2216 ( .A(n3658), .Z(n2934) );
  CANR1X1 U2217 ( .A(n3676), .B(n3675), .C(n3674), .Z(n3677) );
  CIVX1 U2218 ( .A(n3673), .Z(n3675) );
  COR2X1 U2219 ( .A(n3196), .B(n3213), .Z(n2938) );
  COR2X1 U2220 ( .A(n3214), .B(n3213), .Z(n3216) );
  CND3X1 U2221 ( .A(n3219), .B(n3217), .C(n2896), .Z(n3248) );
  CND2X1 U2222 ( .A(n3177), .B(n3102), .Z(n3214) );
  CEOX1 U2223 ( .A(n3665), .B(n3663), .Z(n2972) );
  CNR2X1 U2224 ( .A(n3659), .B(n3020), .Z(n3662) );
  CND3X1 U2225 ( .A(n3303), .B(n2886), .C(n3301), .Z(n3219) );
  CND2IX1 U2226 ( .B(n3189), .A(n2939), .Z(n3110) );
  CNR3X2 U2227 ( .A(n2091), .B(n2089), .C(n2096), .Z(n2165) );
  CIVX1 U2228 ( .A(i[2]), .Z(n2096) );
  CND2IX1 U2229 ( .B(n3209), .A(n2940), .Z(n3210) );
  COR2X1 U2230 ( .A(n3009), .B(n3105), .Z(n3380) );
  CND2X1 U2231 ( .A(n3377), .B(n3104), .Z(n3105) );
  COND1X2 U2232 ( .A(n3303), .B(n3302), .C(n3301), .Z(n3593) );
  CIVX2 U2233 ( .A(n3044), .Z(n3704) );
  CANR1X1 U2234 ( .A(n3666), .B(n3665), .C(n3664), .Z(n3667) );
  CND3XL U2235 ( .A(n2888), .B(n2943), .C(n3202), .Z(n2944) );
  CIVX2 U2236 ( .A(n3322), .Z(n2943) );
  CND2XL U2237 ( .A(n2996), .B(n3712), .Z(n2945) );
  CIVXL U2238 ( .A(n2999), .Z(n2946) );
  COAN1X1 U2239 ( .A(n3414), .B(n3413), .C(n3412), .Z(n2949) );
  CND2X1 U2240 ( .A(n2949), .B(n3411), .Z(n826) );
  CND2XL U2241 ( .A(n3704), .B(n3410), .Z(n3411) );
  COND1XL U2242 ( .A(n3152), .B(n3151), .C(n3150), .Z(n3154) );
  CEOXL U2243 ( .A(opera1[13]), .B(n2879), .Z(n3117) );
  CEOX1 U2244 ( .A(opera1[9]), .B(n2874), .Z(n3131) );
  CEOXL U2245 ( .A(opera1[16]), .B(n2899), .Z(n3174) );
  CND2X1 U2246 ( .A(n2697), .B(n2703), .Z(n2708) );
  CND2X1 U2247 ( .A(n3209), .B(n3195), .Z(n3206) );
  CND2XL U2248 ( .A(n3200), .B(n3194), .Z(n3195) );
  CIVXL U2249 ( .A(res_not_wire[20]), .Z(n2120) );
  CND2IXL U2250 ( .B(n3010), .A(n3145), .Z(n3143) );
  CND2XL U2251 ( .A(n3012), .B(n3130), .Z(n3127) );
  CND2XL U2252 ( .A(n2994), .B(n3126), .Z(n3166) );
  CIVXL U2253 ( .A(c_inop1), .Z(n3151) );
  CND2X1 U2254 ( .A(n2992), .B(n3129), .Z(n3137) );
  CND3XL U2255 ( .A(result[33]), .B(n3154), .C(n3153), .Z(n3743) );
  CIVXL U2256 ( .A(n3153), .Z(n3144) );
  COND2X2 U2257 ( .A(n2942), .B(n3396), .C(n3395), .D(n3394), .Z(n3408) );
  CANR1X2 U2258 ( .A(n3384), .B(n3702), .C(n3383), .Z(n3394) );
  CIVX1 U2259 ( .A(n3221), .Z(n3190) );
  CIVXL U2260 ( .A(n3229), .Z(n3230) );
  CND2X1 U2261 ( .A(n3189), .B(n3188), .Z(n3229) );
  CNR3X2 U2262 ( .A(n2708), .B(n2709), .C(n2715), .Z(n2716) );
  CNR3X2 U2263 ( .A(n2784), .B(n2785), .C(n2791), .Z(n2792) );
  CND2X2 U2264 ( .A(n2773), .B(n2779), .Z(n2784) );
  CIVX2 U2265 ( .A(result[58]), .Z(n2952) );
  CIVXL U2266 ( .A(n3711), .Z(n3714) );
  CND2XL U2267 ( .A(n3696), .B(n3695), .Z(n833) );
  CND2XL U2268 ( .A(n3318), .B(n3317), .Z(n839) );
  CND2XL U2269 ( .A(n3334), .B(n3333), .Z(n836) );
  COND1XL U2270 ( .A(i[20]), .B(n3060), .C(n2211), .Z(n2213) );
  CEOX2 U2271 ( .A(n2921), .B(n2841), .Z(n2840) );
  CND2XL U2272 ( .A(n3763), .B(n2883), .Z(n3369) );
  CIVX2 U2273 ( .A(n2652), .Z(n2954) );
  CNR2IXL U2274 ( .B(result[58]), .A(n3047), .Z(n3243) );
  CNR2XL U2275 ( .A(n2803), .B(n2906), .Z(n2811) );
  CIVX2 U2276 ( .A(n3710), .Z(n2956) );
  CAN2X1 U2277 ( .A(n2954), .B(n2665), .Z(n2957) );
  CAN2XL U2278 ( .A(n2954), .B(n2968), .Z(n2659) );
  CIVX2 U2279 ( .A(n2817), .Z(n2958) );
  CNR2X1 U2280 ( .A(n2906), .B(n2958), .Z(n2959) );
  CNR3X2 U2281 ( .A(n2727), .B(n2728), .C(n2734), .Z(n2735) );
  CNR3X2 U2282 ( .A(n2677), .B(n2671), .C(n2670), .Z(n2678) );
  CNR2XL U2283 ( .A(n3000), .B(n3233), .Z(n2999) );
  CNR2IXL U2284 ( .B(result[58]), .A(n3234), .Z(n3239) );
  CND2X1 U2285 ( .A(n2792), .B(n2798), .Z(n2803) );
  CND2X1 U2286 ( .A(n2986), .B(n3146), .Z(n3099) );
  COR2X1 U2287 ( .A(n3386), .B(n3385), .Z(n3404) );
  CNR2XL U2288 ( .A(n3382), .B(n2083), .Z(n3383) );
  CEOXL U2289 ( .A(n3690), .B(n2961), .Z(n3693) );
  CEOX1 U2290 ( .A(result[36]), .B(n3159), .Z(n3574) );
  CEOX1 U2291 ( .A(n3000), .B(n3233), .Z(n2996) );
  CND2XL U2292 ( .A(n3051), .B(n2783), .Z(n2781) );
  CND2X1 U2293 ( .A(n3309), .B(n3308), .Z(n840) );
  COR2X1 U2294 ( .A(n3018), .B(n3138), .Z(n3621) );
  CANR1XL U2295 ( .A(n3704), .B(n3669), .C(n3668), .Z(n3672) );
  CNR2XL U2296 ( .A(n3025), .B(n3348), .Z(n3351) );
  CIVX1 U2297 ( .A(n3124), .Z(n3130) );
  CND2IXL U2298 ( .B(n3088), .A(n3500), .Z(n3529) );
  CIVXL U2299 ( .A(n3738), .Z(n3739) );
  CEOXL U2300 ( .A(n2960), .B(n2830), .Z(n2835) );
  CEOXL U2301 ( .A(n1983), .B(n1984), .Z(n2960) );
  CND2X1 U2302 ( .A(n2957), .B(n2968), .Z(n2670) );
  CEOXL U2303 ( .A(n2784), .B(n2785), .Z(n2783) );
  CNR2IXL U2304 ( .B(n3323), .A(n3324), .Z(n3325) );
  CND3X1 U2305 ( .A(n3011), .B(n3624), .C(n3623), .Z(n3271) );
  CND2XL U2306 ( .A(n3187), .B(n3186), .Z(n3188) );
  CAOR1X1 U2307 ( .A(n3689), .B(n3688), .C(n3687), .Z(n2961) );
  CND2XL U2308 ( .A(n3377), .B(n3378), .Z(n3379) );
  CND2XL U2309 ( .A(n3189), .B(n3108), .Z(n3109) );
  CNR4X2 U2310 ( .A(n3118), .B(n3119), .C(n3112), .D(n3097), .Z(n3101) );
  CNR2XL U2311 ( .A(n2972), .B(n3044), .Z(n3659) );
  CND2XL U2312 ( .A(n3187), .B(n3184), .Z(n3185) );
  CND2XL U2313 ( .A(n3193), .B(n3183), .Z(n3184) );
  CND2XL U2314 ( .A(n3107), .B(n3103), .Z(n3104) );
  CND2XL U2315 ( .A(n3214), .B(n3213), .Z(n3215) );
  CNR2IXL U2316 ( .B(n3114), .A(n3119), .Z(n3115) );
  CEOXL U2317 ( .A(n3395), .B(n3394), .Z(n3387) );
  CEOXL U2318 ( .A(n2727), .B(n2728), .Z(n2726) );
  CND2XL U2319 ( .A(n3193), .B(n3192), .Z(n3222) );
  CND2XL U2320 ( .A(n3210), .B(n3191), .Z(n3192) );
  CND2XL U2321 ( .A(n3270), .B(n3271), .Z(n3634) );
  CNR2XL U2322 ( .A(n2974), .B(n3044), .Z(n3580) );
  CNR2XL U2323 ( .A(n2975), .B(n3044), .Z(n3604) );
  CNR2XL U2324 ( .A(n2976), .B(n3044), .Z(n3649) );
  CEOXL U2325 ( .A(n3645), .B(n3644), .Z(n2976) );
  CNR2XL U2326 ( .A(n2983), .B(n3044), .Z(n3734) );
  CNR2XL U2327 ( .A(n2984), .B(n3044), .Z(n3751) );
  CNR2XL U2328 ( .A(n2982), .B(n3044), .Z(n3306) );
  CEOXL U2329 ( .A(n3311), .B(n3312), .Z(n2982) );
  CNR2XL U2330 ( .A(n2980), .B(n3044), .Z(n3265) );
  CEOXL U2331 ( .A(n3264), .B(n3263), .Z(n2980) );
  CNR2XL U2332 ( .A(n2981), .B(n3044), .Z(n3281) );
  CEOXL U2333 ( .A(n3632), .B(n3635), .Z(n3636) );
  CNR2IXL U2334 ( .B(n3364), .A(n3044), .Z(n3367) );
  CND2XL U2335 ( .A(n3278), .B(n3279), .Z(n3286) );
  CND2IXL U2336 ( .B(n3247), .A(n3248), .Z(n3712) );
  CNR2XL U2337 ( .A(n2978), .B(n2882), .Z(n3295) );
  CEOXL U2338 ( .A(n3648), .B(n3697), .Z(n2978) );
  CNR2XL U2339 ( .A(n2962), .B(n3044), .Z(n3715) );
  CND2XL U2340 ( .A(n3369), .B(n3068), .Z(n3071) );
  CND2XL U2341 ( .A(n2891), .B(n3069), .Z(n3068) );
  CND2XL U2342 ( .A(n2991), .B(n3135), .Z(n3134) );
  CAN3XL U2343 ( .A(n2881), .B(n3603), .C(n3602), .Z(n2987) );
  CAN3XL U2344 ( .A(n2881), .B(n3639), .C(n3638), .Z(n2988) );
  CAN3XL U2345 ( .A(n2881), .B(n3681), .C(n3680), .Z(n2989) );
  CIVXL U2346 ( .A(n3165), .Z(n3285) );
  CIVX1 U2347 ( .A(n3280), .Z(n3287) );
  CNR3XL U2348 ( .A(n2235), .B(n2885), .C(n100), .Z(n2247) );
  CEOXL U2349 ( .A(n2708), .B(n2709), .Z(n2707) );
  CND2XL U2350 ( .A(n2875), .B(n3535), .Z(n3547) );
  CND2XL U2351 ( .A(n3619), .B(n3620), .Z(n3727) );
  COR2XL U2352 ( .A(n3253), .B(n3750), .Z(n3579) );
  CNR2IXL U2353 ( .B(n2964), .A(n3464), .Z(n3465) );
  CND2IXL U2354 ( .B(n3076), .A(n3500), .Z(n3517) );
  CIVXL U2355 ( .A(n3618), .Z(n3729) );
  CNR2IXL U2356 ( .B(n3743), .A(n3741), .Z(n3366) );
  CIVX1 U2357 ( .A(n2830), .Z(n1982) );
  CEOXL U2358 ( .A(opera2[5]), .B(n1983), .Z(n2677) );
  CND2XL U2359 ( .A(n3051), .B(n2821), .Z(n2819) );
  CND2XL U2360 ( .A(n2881), .B(n3477), .Z(n3480) );
  CND2XL U2361 ( .A(n3051), .B(n2816), .Z(n2814) );
  CND2XL U2362 ( .A(n2881), .B(n3560), .Z(n3563) );
  CND2XL U2363 ( .A(n2809), .B(n3050), .Z(n2807) );
  CND2XL U2364 ( .A(n2881), .B(n3555), .Z(n3558) );
  CND2XL U2365 ( .A(n2790), .B(n3050), .Z(n2788) );
  CEOXL U2366 ( .A(opera2[8]), .B(n1983), .Z(n2696) );
  CND2XL U2367 ( .A(n2881), .B(n3459), .Z(n3462) );
  CND2XL U2368 ( .A(n3051), .B(n2778), .Z(n2776) );
  CND2XL U2369 ( .A(n2881), .B(n3542), .Z(n3545) );
  CNR2IXL U2370 ( .B(result[49]), .A(n3752), .Z(n3316) );
  CEOXL U2371 ( .A(opera2[11]), .B(n1983), .Z(n2715) );
  CND2XL U2372 ( .A(n3704), .B(n3703), .Z(n3707) );
  CND2XL U2373 ( .A(n2881), .B(n3710), .Z(n3249) );
  CND3X2 U2374 ( .A(i[28]), .B(n2000), .C(i[29]), .Z(n2233) );
  CND2XL U2375 ( .A(n3051), .B(n2764), .Z(n2762) );
  CND2XL U2376 ( .A(n2881), .B(n3536), .Z(n3539) );
  CND2XL U2377 ( .A(n3051), .B(n2759), .Z(n2757) );
  CNR2IXL U2378 ( .B(result[54]), .A(n3046), .Z(n3349) );
  CNR2IXL U2379 ( .B(result[52]), .A(n3752), .Z(n3332) );
  CNR2XL U2380 ( .A(n3734), .B(n3021), .Z(n3737) );
  CND2XL U2381 ( .A(n3737), .B(n3736), .Z(n850) );
  CNR2XL U2382 ( .A(n3022), .B(n3265), .Z(n3268) );
  CND2XL U2383 ( .A(n3268), .B(n3267), .Z(n852) );
  CND2XL U2384 ( .A(n3590), .B(n3589), .Z(n854) );
  CENXL U2385 ( .A(n3585), .B(n3584), .Z(n3587) );
  CND2XL U2386 ( .A(n3631), .B(n3630), .Z(n849) );
  CND2XL U2387 ( .A(n3299), .B(n3298), .Z(n843) );
  CAN3XL U2388 ( .A(n2881), .B(n3731), .C(n3262), .Z(n3022) );
  CAN3XL U2389 ( .A(n2881), .B(n3733), .C(n3732), .Z(n3021) );
  CND2XL U2390 ( .A(n3690), .B(n3221), .Z(n3232) );
  COND1X1 U2391 ( .A(n3232), .B(n2894), .C(n3231), .Z(n3247) );
  CEOXL U2392 ( .A(opera1[17]), .B(n2899), .Z(n3213) );
  CND2XL U2393 ( .A(i[4]), .B(n2169), .Z(n2175) );
  CND2XL U2394 ( .A(i[6]), .B(n2178), .Z(n2177) );
  CND2XL U2395 ( .A(i[1]), .B(n2173), .Z(n2172) );
  CEOXL U2396 ( .A(opera2[17]), .B(n1983), .Z(n2753) );
  COND11XL U2397 ( .A(n3060), .B(i[12]), .C(n2191), .D(n2192), .Z(n942) );
  COND11XL U2398 ( .A(n3060), .B(i[26]), .C(n2223), .D(n2224), .Z(n928) );
  COND11XL U2399 ( .A(n3060), .B(i[8]), .C(n2181), .D(n2182), .Z(n946) );
  CEOXL U2400 ( .A(opera1[18]), .B(n2899), .Z(n3196) );
  CEOXL U2401 ( .A(opera2[14]), .B(n1983), .Z(n2734) );
  CEOXL U2402 ( .A(n3710), .B(n108), .Z(n3716) );
  CND2XL U2403 ( .A(res_not_wire[28]), .B(n3476), .Z(n3564) );
  CANR2XL U2404 ( .A(result[34]), .B(n3057), .C(n3053), .D(n3760), .Z(n2285)
         );
  CANR2XL U2405 ( .A(result[35]), .B(n3055), .C(n3053), .D(n2046), .Z(n2286)
         );
  CANR2XL U2406 ( .A(result[32]), .B(n3057), .C(n3053), .D(n2099), .Z(n2283)
         );
  CANR2XL U2407 ( .A(result[37]), .B(n3055), .C(n3053), .D(n3002), .Z(n2288)
         );
  CNR2IXL U2408 ( .B(result[33]), .A(n3369), .Z(n3372) );
  CEOXL U2409 ( .A(n3482), .B(n134), .Z(n3080) );
  CND2XL U2410 ( .A(n3704), .B(n3387), .Z(n3390) );
  CND2XL U2411 ( .A(n2881), .B(n3421), .Z(n3424) );
  CND2XL U2412 ( .A(n2881), .B(n3434), .Z(n3437) );
  CND2XL U2413 ( .A(n2881), .B(n3487), .Z(n3490) );
  CND2XL U2414 ( .A(n2881), .B(n3492), .Z(n3495) );
  CND2XL U2415 ( .A(n2881), .B(n3501), .Z(n3504) );
  CND2XL U2416 ( .A(n2881), .B(n3506), .Z(n3509) );
  CND2XL U2417 ( .A(n2881), .B(n3518), .Z(n3521) );
  CND2XL U2418 ( .A(n2881), .B(n3524), .Z(n3527) );
  CND2XL U2419 ( .A(n2714), .B(n3050), .Z(n2712) );
  COND4CXL U2420 ( .A(n2161), .B(n2154), .C(n2169), .D(i[5]), .Z(n2168) );
  CNR2XL U2421 ( .A(n2997), .B(n2882), .Z(n3586) );
  CEOXL U2422 ( .A(res_not_wire[34]), .B(n3750), .Z(n2997) );
  CNR2XL U2423 ( .A(n2998), .B(n2882), .Z(n3627) );
  CNR2XL U2424 ( .A(n3007), .B(n2882), .Z(n3668) );
  CEOXL U2425 ( .A(n114), .B(n2934), .Z(n3007) );
  CNR2IXL U2426 ( .B(result[31]), .A(n3752), .Z(n3079) );
  CNR2IXL U2427 ( .B(result[43]), .A(n3045), .Z(n3292) );
  CNR2IXL U2428 ( .B(result[45]), .A(n3752), .Z(n3297) );
  CNR2IXL U2429 ( .B(result[60]), .A(n3045), .Z(n3388) );
  CAN2X1 U2430 ( .A(n2965), .B(res_not_wire[16]), .Z(n2964) );
  COR2XL U2431 ( .A(n3006), .B(n3142), .Z(n3619) );
  CND2XL U2432 ( .A(n2881), .B(n3446), .Z(n3449) );
  CANR2XL U2433 ( .A(n3704), .B(n3273), .C(n2881), .D(n3272), .Z(n3276) );
  CANR2XL U2434 ( .A(n3704), .B(n3291), .C(n2881), .D(n3290), .Z(n3294) );
  CNR2XL U2435 ( .A(n3649), .B(n3019), .Z(n3652) );
  CND2XL U2436 ( .A(n3652), .B(n3651), .Z(n844) );
  CNR2XL U2437 ( .A(n3023), .B(n3281), .Z(n3284) );
  CND2XL U2438 ( .A(n3284), .B(n3283), .Z(n846) );
  CND2XL U2439 ( .A(n3719), .B(n3718), .Z(n831) );
  COND4CXL U2440 ( .A(n2161), .B(n2153), .C(n2178), .D(i[7]), .Z(n2179) );
  CAN3XL U2441 ( .A(n2881), .B(n3646), .C(n3277), .Z(n3023) );
  CAN3XL U2442 ( .A(n2881), .B(n3656), .C(n3300), .Z(n3024) );
  CAN3XL U2443 ( .A(n2881), .B(n3336), .C(n3335), .Z(n3025) );
  CAN3XL U2444 ( .A(n2881), .B(n3648), .C(n3647), .Z(n3019) );
  CAN3XL U2445 ( .A(n2881), .B(n3658), .C(n3657), .Z(n3020) );
  CNR2IXL U2446 ( .B(res_not_wire[18]), .A(n3058), .Z(n3355) );
  CNR2IXL U2447 ( .B(res_not_wire[12]), .A(n3058), .Z(n3361) );
  CNR2IXL U2448 ( .B(res_not_wire[36]), .A(n3058), .Z(n3721) );
  CMXI2XL U2449 ( .A0(n3052), .A1(n3057), .S(result[36]), .Z(n3720) );
  CNR2IXL U2450 ( .B(res_not_wire[24]), .A(n3058), .Z(n3722) );
  CMXI2XL U2451 ( .A0(n3052), .A1(n3057), .S(result[33]), .Z(n3723) );
  CEOXL U2452 ( .A(n3476), .B(res_not_wire[28]), .Z(n3477) );
  CEOXL U2453 ( .A(opera2[20]), .B(n1983), .Z(n2772) );
  CENX1 U2454 ( .A(n2966), .B(n3559), .Z(n3560) );
  CND2XL U2455 ( .A(n3553), .B(n3470), .Z(n3559) );
  CNR2IXL U2456 ( .B(res_not_wire[26]), .A(n3554), .Z(n3470) );
  COR2XL U2457 ( .A(n3028), .B(n3087), .Z(n3254) );
  CND2IXL U2458 ( .B(n142), .A(n3001), .Z(n3258) );
  CIVXL U2459 ( .A(i[4]), .Z(n2154) );
  CIVXL U2460 ( .A(i[3]), .Z(n2148) );
  CEOXL U2461 ( .A(opera2[23]), .B(n1983), .Z(n2791) );
  CNR2IXL U2462 ( .B(res_not_wire[16]), .A(n3258), .Z(n3259) );
  CND2IXL U2463 ( .B(res_not_wire[12]), .A(n3512), .Z(n3438) );
  CND2IXL U2464 ( .B(res_not_wire[18]), .A(n3531), .Z(n3450) );
  CIVXL U2465 ( .A(res_not_wire[32]), .Z(n3370) );
  CEOXL U2466 ( .A(opera2[26]), .B(n1983), .Z(n2810) );
  CEOXL U2467 ( .A(opera2[29]), .B(n1983), .Z(n2829) );
  CEOXL U2468 ( .A(res_not_wire[4]), .B(n3034), .Z(n3421) );
  CEOXL U2469 ( .A(n3486), .B(n164), .Z(n3487) );
  CIVXL U2470 ( .A(result[32]), .Z(n2099) );
  CIVXL U2471 ( .A(result[34]), .Z(n3760) );
  CIVX2 U2472 ( .A(n3049), .Z(n3048) );
  CIVX2 U2473 ( .A(n3049), .Z(n3047) );
  CIVX2 U2474 ( .A(n3049), .Z(n3046) );
  CIVX2 U2475 ( .A(n3049), .Z(n3045) );
  CIVX2 U2476 ( .A(n3060), .Z(n3059) );
  CIVX2 U2477 ( .A(n2885), .Z(n3058) );
  CIVX2 U2478 ( .A(n3369), .Z(n3754) );
  CNIVX1 U2479 ( .A(n2246), .Z(n3055) );
  COND1XL U2480 ( .A(n2889), .B(n3180), .C(n3179), .Z(n3181) );
  CND2X1 U2481 ( .A(n2885), .B(n2236), .Z(n2170) );
  CNIVX1 U2482 ( .A(n2246), .Z(n3056) );
  CNIVX1 U2483 ( .A(n2246), .Z(n3057) );
  CND3XL U2484 ( .A(n3123), .B(n2985), .C(n3139), .Z(n3124) );
  CND2X1 U2485 ( .A(n3180), .B(n2889), .Z(n3179) );
  CND2X1 U2486 ( .A(n2888), .B(n3202), .Z(n3327) );
  COND1XL U2487 ( .A(n2087), .B(n3060), .C(n2170), .Z(n2178) );
  COND1XL U2488 ( .A(n2088), .B(n3060), .C(n2170), .Z(n2169) );
  COND1XL U2489 ( .A(n2001), .B(n3060), .C(n2170), .Z(n2225) );
  COND1XL U2490 ( .A(n2010), .B(n3060), .C(n2170), .Z(n2188) );
  COND1XL U2491 ( .A(n2007), .B(n3060), .C(n2170), .Z(n2206) );
  CNIVX1 U2492 ( .A(n2247), .Z(n3054) );
  CNIVX1 U2493 ( .A(n2247), .Z(n3053) );
  CNIVX1 U2494 ( .A(n2247), .Z(n3052) );
  CAN2X1 U2495 ( .A(n3624), .B(n3623), .Z(n3625) );
  CAN2X1 U2496 ( .A(n2236), .B(n2101), .Z(n2238) );
  CNR2IX1 U2497 ( .B(n3278), .A(n3285), .Z(n3171) );
  CANR1XL U2498 ( .A(n3117), .B(n3167), .C(n2889), .Z(n3173) );
  CANR3X1 U2499 ( .A(n3338), .B(n3599), .C(n3224), .D(n3312), .Z(n3339) );
  CANR1XL U2500 ( .A(n3131), .B(n3134), .C(n3130), .Z(n3132) );
  CNR3X2 U2501 ( .A(n2829), .B(n2823), .C(n2822), .Z(n2830) );
  CANR1XL U2502 ( .A(n2209), .B(n3059), .C(n1989), .Z(n2211) );
  CNR3X2 U2503 ( .A(n2753), .B(n2747), .C(n2746), .Z(n2754) );
  CNR2X1 U2504 ( .A(n2977), .B(n3044), .Z(n3682) );
  CEOX1 U2505 ( .A(n3014), .B(n3677), .Z(n2977) );
  COND1XL U2506 ( .A(n3135), .B(n2991), .C(n3134), .Z(n3136) );
  CANR1XL U2507 ( .A(n2091), .B(n3059), .C(n2173), .Z(n2162) );
  CND3XL U2508 ( .A(n3301), .B(n3302), .C(n2886), .Z(n3218) );
  CND2X1 U2509 ( .A(n2846), .B(n3768), .Z(n2236) );
  CNR2X1 U2510 ( .A(n2979), .B(n3044), .Z(n3348) );
  CEOX1 U2511 ( .A(n3689), .B(n3347), .Z(n2979) );
  CEOX1 U2512 ( .A(n3286), .B(n3280), .Z(n2981) );
  CND2X1 U2513 ( .A(n3059), .B(n2215), .Z(n2201) );
  CND2X1 U2514 ( .A(n3379), .B(n3386), .Z(n3382) );
  COR2X1 U2515 ( .A(n3210), .B(n3191), .Z(n3193) );
  COR2X1 U2516 ( .A(n3193), .B(n3183), .Z(n3187) );
  COR2X1 U2517 ( .A(n3187), .B(n3186), .Z(n3189) );
  COR2X1 U2518 ( .A(n3110), .B(n3106), .Z(n3107) );
  COR2X1 U2519 ( .A(n3107), .B(n3103), .Z(n3377) );
  CNR2X1 U2520 ( .A(n2996), .B(n2999), .Z(n3235) );
  CEOX1 U2521 ( .A(n3729), .B(n3728), .Z(n2983) );
  CENX1 U2522 ( .A(n3745), .B(n3744), .Z(n2984) );
  CNR2IX1 U2523 ( .B(n3320), .A(n3044), .Z(n3331) );
  CND2X1 U2524 ( .A(n3127), .B(n3125), .Z(n3133) );
  CND2X1 U2525 ( .A(n3010), .B(n3139), .Z(n3160) );
  COR2X1 U2526 ( .A(n3199), .B(n3198), .Z(n3200) );
  CND3XL U2527 ( .A(n3375), .B(n3374), .C(n3373), .Z(n856) );
  CNR2X1 U2528 ( .A(n3372), .B(n2897), .Z(n3373) );
  CND2X1 U2529 ( .A(n3014), .B(n3674), .Z(n3342) );
  CND2X1 U2530 ( .A(n2240), .B(n3062), .Z(n3063) );
  CND2X1 U2531 ( .A(n3686), .B(n3337), .Z(n3221) );
  CND2X1 U2532 ( .A(n3101), .B(n3100), .Z(n3175) );
  CND2X1 U2533 ( .A(n3204), .B(n3653), .Z(n3205) );
  COR2X1 U2534 ( .A(n2938), .B(n3214), .Z(n3199) );
  CND2X1 U2535 ( .A(n3621), .B(n3618), .Z(n3624) );
  CIVX2 U2536 ( .A(n3392), .Z(n3402) );
  CIVX2 U2537 ( .A(n2171), .Z(n2088) );
  CND2X1 U2538 ( .A(n3227), .B(n3228), .Z(n3674) );
  CND2X1 U2539 ( .A(n3676), .B(n3226), .Z(n3227) );
  CIVX2 U2540 ( .A(n2223), .Z(n2001) );
  CIVX2 U2541 ( .A(n2186), .Z(n2010) );
  CND2IX1 U2542 ( .B(n2999), .A(n3248), .Z(n3237) );
  CAN2X1 U2543 ( .A(n3148), .B(n3017), .Z(n2986) );
  CANR1XL U2544 ( .A(n3633), .B(n3269), .C(n3632), .Z(n3163) );
  CND3X1 U2545 ( .A(n3633), .B(n3270), .C(n3271), .Z(n3162) );
  CAN3X2 U2546 ( .A(n2881), .B(n3750), .C(n3749), .Z(n2990) );
  CIVX2 U2547 ( .A(n2232), .Z(n2000) );
  CIVX2 U2548 ( .A(n3417), .Z(n3491) );
  CIVX2 U2549 ( .A(n2176), .Z(n2087) );
  CANR1XL U2550 ( .A(n2232), .B(n3059), .C(n1989), .Z(n2228) );
  CANR1XL U2551 ( .A(n2842), .B(n3758), .C(n2244), .Z(n3062) );
  CNR3XL U2552 ( .A(n3531), .B(n3258), .C(n3254), .Z(n3476) );
  CND2X1 U2553 ( .A(n3764), .B(n2102), .Z(n2242) );
  COND1XL U2554 ( .A(n2215), .B(n3060), .C(n2170), .Z(n2202) );
  COND2X1 U2555 ( .A(n2228), .B(n2093), .C(n3060), .D(n2229), .Z(n926) );
  CENX1 U2556 ( .A(n2995), .B(n3288), .Z(n3291) );
  CANR1XL U2557 ( .A(n3287), .B(n3286), .C(n3285), .Z(n3288) );
  CANR1XL U2558 ( .A(n3729), .B(n3727), .C(n3622), .Z(n3626) );
  CENX1 U2559 ( .A(n3731), .B(n3612), .Z(n3613) );
  CNR3XL U2560 ( .A(n3364), .B(n2235), .C(n3763), .Z(n3368) );
  CENX1 U2561 ( .A(opera1[14]), .B(n2873), .Z(n3176) );
  CENX1 U2562 ( .A(res_not_wire[52]), .B(n2935), .Z(n3329) );
  CEOX1 U2563 ( .A(opera2[3]), .B(opera2_63), .Z(n2665) );
  CENX1 U2564 ( .A(res_not_wire[58]), .B(n3016), .Z(n3246) );
  CANR1XL U2565 ( .A(result[59]), .B(n3754), .C(n3243), .Z(n3244) );
  CND3XL U2566 ( .A(n3381), .B(n3704), .C(n3242), .Z(n3245) );
  CEOX1 U2567 ( .A(result[49]), .B(n3223), .Z(n3312) );
  CEOX1 U2568 ( .A(result[42]), .B(n3133), .Z(n3632) );
  COND1XL U2569 ( .A(n3182), .B(result[47]), .C(n3304), .Z(n3592) );
  CENX1 U2570 ( .A(n2878), .B(opera1[0]), .Z(n3152) );
  CANR2X1 U2571 ( .A(result[9]), .B(n3055), .C(n3052), .D(n2059), .Z(n2260) );
  CANR2X1 U2572 ( .A(result[7]), .B(n3055), .C(n3052), .D(n2060), .Z(n2258) );
  COND11X1 U2573 ( .A(n2201), .B(i[23]), .C(n2003), .D(n2216), .Z(n931) );
  COND11X1 U2574 ( .A(n2212), .B(i[22]), .C(n2147), .D(n2214), .Z(n932) );
  CND2X1 U2575 ( .A(i[8]), .B(n2183), .Z(n2182) );
  COND11X1 U2576 ( .A(n2201), .B(i[17]), .C(n2149), .D(n2203), .Z(n937) );
  CANR2X1 U2577 ( .A(result[19]), .B(n3056), .C(n3053), .D(n2054), .Z(n2270)
         );
  CEOX1 U2578 ( .A(result[50]), .B(n3203), .Z(n3322) );
  CENX1 U2579 ( .A(result[35]), .B(n2970), .Z(n3584) );
  CENX1 U2580 ( .A(result[45]), .B(n3173), .Z(n3644) );
  COND1XL U2581 ( .A(n3132), .B(result[41]), .C(n3633), .Z(n3269) );
  CND2X1 U2582 ( .A(result[56]), .B(n3230), .Z(n3231) );
  COND2X1 U2583 ( .A(n1986), .B(n2149), .C(i[16]), .D(n2201), .Z(n938) );
  CANR1XL U2584 ( .A(result[60]), .B(n3754), .C(n3705), .Z(n3706) );
  CANR1XL U2585 ( .A(result[62]), .B(n3754), .C(n3397), .Z(n3398) );
  CND2X1 U2586 ( .A(n3051), .B(n2914), .Z(n2641) );
  CANR1XL U2587 ( .A(result[63]), .B(n3754), .C(n3403), .Z(n3412) );
  CND2X1 U2588 ( .A(result[41]), .B(n3132), .Z(n3633) );
  CND4X1 U2589 ( .A(res_not_wire[26]), .B(n3553), .C(res_not_wire[24]), .D(
        n3078), .Z(n3087) );
  COND1XL U2590 ( .A(n3405), .B(result[62]), .C(n3029), .Z(n3406) );
  CANR1X1 U2591 ( .A(n2941), .B(n3408), .C(n3407), .Z(n3409) );
  CND3XL U2592 ( .A(n2881), .B(n3482), .C(n3481), .Z(n3485) );
  CND2X1 U2593 ( .A(n2657), .B(n3050), .Z(n2655) );
  CND2X1 U2594 ( .A(result[47]), .B(n3182), .Z(n3304) );
  CEOX1 U2595 ( .A(result[44]), .B(n2969), .Z(n2995) );
  COND1XL U2596 ( .A(n2882), .B(n3573), .C(n3572), .Z(n919) );
  CNR2X1 U2597 ( .A(n3253), .B(n132), .Z(n3089) );
  CNR2IX1 U2598 ( .B(result[4]), .A(n3045), .Z(n3422) );
  CNR2IX1 U2599 ( .B(result[6]), .A(n3047), .Z(n3427) );
  CNR2IX1 U2600 ( .B(result[8]), .A(n3048), .Z(n3431) );
  CNR2IX1 U2601 ( .B(result[10]), .A(n3046), .Z(n3435) );
  CNR2IX1 U2602 ( .B(result[12]), .A(n3047), .Z(n3439) );
  CNR2IX1 U2603 ( .B(result[14]), .A(n3045), .Z(n3443) );
  CNR2IX1 U2604 ( .B(result[16]), .A(n3046), .Z(n3447) );
  CNR2IX1 U2605 ( .B(result[20]), .A(n3048), .Z(n3456) );
  CNR2IX1 U2606 ( .B(result[22]), .A(n3046), .Z(n3460) );
  CNR2IX1 U2607 ( .B(result[24]), .A(n3047), .Z(n3467) );
  CNR2IX1 U2608 ( .B(result[26]), .A(n3048), .Z(n3473) );
  CNR2IX1 U2609 ( .B(result[28]), .A(n3045), .Z(n3478) );
  CNR2IX1 U2610 ( .B(result[1]), .A(n3048), .Z(n3488) );
  CNR2IX1 U2611 ( .B(result[3]), .A(n3045), .Z(n3493) );
  CNR2IX1 U2612 ( .B(result[5]), .A(n3048), .Z(n3497) );
  CNR2IX1 U2613 ( .B(result[7]), .A(n3046), .Z(n3502) );
  CNR2IX1 U2614 ( .B(result[9]), .A(n3046), .Z(n3507) );
  CNR2IX1 U2615 ( .B(result[11]), .A(n3047), .Z(n3513) );
  CNR2IX1 U2616 ( .B(result[13]), .A(n3045), .Z(n3519) );
  CNR2IX1 U2617 ( .B(result[15]), .A(n3045), .Z(n3525) );
  CNR2IX1 U2618 ( .B(result[17]), .A(n3046), .Z(n3532) );
  CNR2IX1 U2619 ( .B(result[19]), .A(n3047), .Z(n3537) );
  CNR2IX1 U2620 ( .B(result[21]), .A(n3045), .Z(n3543) );
  CNR2IX1 U2621 ( .B(result[23]), .A(n3046), .Z(n3550) );
  CNR2IX1 U2622 ( .B(result[25]), .A(n3048), .Z(n3556) );
  COND1XL U2623 ( .A(n140), .B(n3058), .C(n2276), .Z(n894) );
  CANR2X1 U2624 ( .A(result[25]), .B(n3055), .C(n3053), .D(n2051), .Z(n2276)
         );
  COND1XL U2625 ( .A(n138), .B(n3058), .C(n2278), .Z(n892) );
  CANR2X1 U2626 ( .A(result[27]), .B(n3057), .C(n3053), .D(n2050), .Z(n2278)
         );
  COND1XL U2627 ( .A(n136), .B(n3058), .C(n2280), .Z(n890) );
  CANR2X1 U2628 ( .A(result[29]), .B(n3056), .C(n3053), .D(n2049), .Z(n2280)
         );
  COND1XL U2629 ( .A(n124), .B(n3058), .C(n2292), .Z(n878) );
  CANR2X1 U2630 ( .A(result[41]), .B(n3057), .C(n3054), .D(n2035), .Z(n2292)
         );
  COND1XL U2631 ( .A(n114), .B(n3058), .C(n2302), .Z(n868) );
  CANR2X1 U2632 ( .A(result[51]), .B(n3057), .C(n3054), .D(n3008), .Z(n2302)
         );
  COND1XL U2633 ( .A(n3058), .B(n2106), .C(n2848), .Z(n793) );
  CANR2X1 U2634 ( .A(result[63]), .B(n3057), .C(n3054), .D(n3769), .Z(n2848)
         );
  COND1XL U2635 ( .A(n152), .B(n3058), .C(n2264), .Z(n906) );
  CANR2X1 U2636 ( .A(result[13]), .B(n3056), .C(n3052), .D(n2057), .Z(n2264)
         );
  COND1XL U2637 ( .A(n150), .B(n3058), .C(n2266), .Z(n904) );
  CANR2X1 U2638 ( .A(result[15]), .B(n3056), .C(n3054), .D(n2056), .Z(n2266)
         );
  COND1XL U2639 ( .A(n148), .B(n3058), .C(n2268), .Z(n902) );
  CANR2X1 U2640 ( .A(result[17]), .B(n3056), .C(n3054), .D(n2055), .Z(n2268)
         );
  COND1XL U2641 ( .A(n3058), .B(n3761), .C(n2311), .Z(n859) );
  CANR2X1 U2642 ( .A(result[60]), .B(n3057), .C(n3053), .D(n2083), .Z(n2311)
         );
  COND1XL U2643 ( .A(n112), .B(n3058), .C(n2304), .Z(n866) );
  CANR2X1 U2644 ( .A(result[53]), .B(n3057), .C(n3054), .D(n3003), .Z(n2304)
         );
  COND1XL U2645 ( .A(n130), .B(n3058), .C(n2286), .Z(n884) );
  CANR2X1 U2646 ( .A(result[23]), .B(n3056), .C(n3052), .D(n2052), .Z(n2274)
         );
  COND1XL U2647 ( .A(n116), .B(n3058), .C(n2300), .Z(n870) );
  CANR2X1 U2648 ( .A(result[49]), .B(n3057), .C(n3054), .D(n2137), .Z(n2300)
         );
  COND1XL U2649 ( .A(n118), .B(n3058), .C(n2298), .Z(n872) );
  CANR2X1 U2650 ( .A(result[47]), .B(n3057), .C(n3054), .D(n3759), .Z(n2298)
         );
  COND1XL U2651 ( .A(n110), .B(n3058), .C(n2306), .Z(n864) );
  CANR2X1 U2652 ( .A(result[55]), .B(n3057), .C(n3054), .D(n3004), .Z(n2306)
         );
  COND1XL U2653 ( .A(n108), .B(n3058), .C(n2308), .Z(n862) );
  CANR2X1 U2654 ( .A(result[57]), .B(n3057), .C(n3052), .D(n3000), .Z(n2308)
         );
  COND1XL U2655 ( .A(n3058), .B(n2024), .C(n2310), .Z(n860) );
  CANR2X1 U2656 ( .A(result[59]), .B(n3057), .C(n3053), .D(n3009), .Z(n2310)
         );
  COND1XL U2657 ( .A(n3058), .B(n3546), .C(n2273), .Z(n897) );
  CANR2X1 U2658 ( .A(result[22]), .B(n3056), .C(n3053), .D(n2068), .Z(n2273)
         );
  COND1XL U2659 ( .A(n144), .B(n3058), .C(n2272), .Z(n898) );
  CANR2X1 U2660 ( .A(result[21]), .B(n3056), .C(n3054), .D(n2053), .Z(n2272)
         );
  COND1XL U2661 ( .A(n3058), .B(n2020), .C(n2312), .Z(n858) );
  CANR2X1 U2662 ( .A(result[61]), .B(n3057), .C(n3052), .D(n2942), .Z(n2312)
         );
  COND1XL U2663 ( .A(n3058), .B(n3370), .C(n2283), .Z(n887) );
  COND1XL U2664 ( .A(n3058), .B(n2018), .C(n2313), .Z(n857) );
  CANR2X1 U2665 ( .A(result[62]), .B(n3057), .C(n3052), .D(n3762), .Z(n2313)
         );
  COND1XL U2666 ( .A(n128), .B(n3058), .C(n2288), .Z(n882) );
  COND1XL U2667 ( .A(n3058), .B(n3084), .C(n2307), .Z(n863) );
  CANR2X1 U2668 ( .A(result[56]), .B(n3057), .C(n3054), .D(n2144), .Z(n2307)
         );
  COND1XL U2669 ( .A(n3058), .B(n2013), .C(n2309), .Z(n861) );
  CANR2X1 U2670 ( .A(result[58]), .B(n3057), .C(n3054), .D(n2952), .Z(n2309)
         );
  COND1XL U2671 ( .A(n160), .B(n3058), .C(n2256), .Z(n914) );
  CANR2X1 U2672 ( .A(result[5]), .B(n3055), .C(n3052), .D(n2061), .Z(n2256) );
  COND1XL U2673 ( .A(n164), .B(n3058), .C(n2252), .Z(n918) );
  CANR2X1 U2674 ( .A(result[1]), .B(n3055), .C(n3052), .D(n2063), .Z(n2252) );
  COND1XL U2675 ( .A(n154), .B(n3058), .C(n2262), .Z(n908) );
  CANR2X1 U2676 ( .A(result[11]), .B(n3055), .C(n3052), .D(n2058), .Z(n2262)
         );
  COND1XL U2677 ( .A(n162), .B(n3058), .C(n2254), .Z(n916) );
  CANR2X1 U2678 ( .A(result[3]), .B(n3055), .C(n3052), .D(n2062), .Z(n2254) );
  COND1XL U2679 ( .A(n3058), .B(n3767), .C(n2281), .Z(n889) );
  CANR2X1 U2680 ( .A(result[30]), .B(n3055), .C(n3053), .D(n2064), .Z(n2281)
         );
  COND1XL U2681 ( .A(n3058), .B(n3471), .C(n2277), .Z(n893) );
  CANR2X1 U2682 ( .A(result[26]), .B(n3057), .C(n3053), .D(n2066), .Z(n2277)
         );
  COND1XL U2683 ( .A(n3058), .B(n2131), .C(n2279), .Z(n891) );
  CANR2X1 U2684 ( .A(result[28]), .B(n3055), .C(n3053), .D(n2065), .Z(n2279)
         );
  COND1XL U2685 ( .A(n3058), .B(n3577), .C(n2285), .Z(n885) );
  COND1XL U2686 ( .A(n3058), .B(n2128), .C(n2297), .Z(n873) );
  CANR2X1 U2687 ( .A(result[46]), .B(n3057), .C(n3054), .D(n3026), .Z(n2297)
         );
  COND1XL U2688 ( .A(n3058), .B(n3766), .C(n2299), .Z(n871) );
  CANR2X1 U2689 ( .A(result[48]), .B(n3057), .C(n3054), .D(n2138), .Z(n2299)
         );
  COND1XL U2690 ( .A(n3058), .B(n3655), .C(n2301), .Z(n869) );
  CANR2X1 U2691 ( .A(result[50]), .B(n3057), .C(n3054), .D(n3005), .Z(n2301)
         );
  COND1XL U2692 ( .A(n3058), .B(n2125), .C(n2303), .Z(n867) );
  CANR2X1 U2693 ( .A(result[52]), .B(n3057), .C(n3054), .D(n2136), .Z(n2303)
         );
  COND1XL U2694 ( .A(n3058), .B(n3765), .C(n2305), .Z(n865) );
  CANR2X1 U2695 ( .A(result[54]), .B(n3057), .C(n3054), .D(n2135), .Z(n2305)
         );
  COND1XL U2696 ( .A(n3058), .B(n3036), .C(n2265), .Z(n905) );
  CANR2X1 U2697 ( .A(result[14]), .B(n3056), .C(n3052), .D(n2072), .Z(n2265)
         );
  COND1XL U2698 ( .A(n3058), .B(n2120), .C(n2271), .Z(n899) );
  CANR2X1 U2699 ( .A(result[20]), .B(n3056), .C(n3054), .D(n2069), .Z(n2271)
         );
  COND1XL U2700 ( .A(n3058), .B(n3528), .C(n2267), .Z(n903) );
  CANR2X1 U2701 ( .A(result[16]), .B(n3056), .C(n3053), .D(n2071), .Z(n2267)
         );
  COND1XL U2702 ( .A(n3058), .B(n3352), .C(n2245), .Z(n920) );
  CANR2X1 U2703 ( .A(result[0]), .B(n3055), .C(n3052), .D(n3763), .Z(n2245) );
  COND1XL U2704 ( .A(n3058), .B(n2123), .C(n2259), .Z(n911) );
  CANR2X1 U2705 ( .A(result[8]), .B(n3055), .C(n3052), .D(n2075), .Z(n2259) );
  COND1XL U2706 ( .A(n3058), .B(n3415), .C(n2253), .Z(n917) );
  CANR2X1 U2707 ( .A(result[2]), .B(n3055), .C(n3052), .D(n2078), .Z(n2253) );
  COND1XL U2708 ( .A(n3058), .B(n2116), .C(n2261), .Z(n909) );
  CANR2X1 U2709 ( .A(result[10]), .B(n3055), .C(n3052), .D(n2074), .Z(n2261)
         );
  COND4CX1 U2710 ( .A(n2228), .B(n2230), .C(n2094), .D(n2231), .Z(n925) );
  CNIVX4 U2711 ( .A(n3746), .Z(n3044) );
  CAN2X1 U2712 ( .A(res_not_wire[18]), .B(n2875), .Z(n3001) );
  COND1XL U2713 ( .A(n3058), .B(n2118), .C(n2255), .Z(n915) );
  CANR2X1 U2714 ( .A(result[4]), .B(n3055), .C(n3052), .D(n2077), .Z(n2255) );
  COR2X1 U2715 ( .A(n3003), .B(n3211), .Z(n3228) );
  CND2X1 U2716 ( .A(n2148), .B(n2154), .Z(n2849) );
  COR2X1 U2717 ( .A(n3005), .B(n3203), .Z(n3653) );
  CND2X1 U2718 ( .A(n3228), .B(n3212), .Z(n3224) );
  CNR2IX1 U2719 ( .B(result[62]), .A(n3046), .Z(n3403) );
  COR2X1 U2720 ( .A(n3008), .B(n3201), .Z(n3204) );
  CNR2IX1 U2721 ( .B(n2903), .A(n3084), .Z(n3096) );
  CND3XL U2722 ( .A(n3391), .B(n3390), .C(n3389), .Z(n828) );
  CANR1XL U2723 ( .A(result[61]), .B(n3754), .C(n3388), .Z(n3389) );
  CND3XL U2724 ( .A(n2667), .B(n3424), .C(n3423), .Z(n821) );
  CANR1XL U2725 ( .A(result[5]), .B(n2891), .C(n3422), .Z(n3423) );
  CND3XL U2726 ( .A(n2681), .B(n3429), .C(n3428), .Z(n819) );
  CANR1XL U2727 ( .A(result[7]), .B(n2891), .C(n3427), .Z(n3428) );
  CND3XL U2728 ( .A(n2705), .B(n3437), .C(n3436), .Z(n815) );
  CANR1XL U2729 ( .A(result[11]), .B(n2891), .C(n3435), .Z(n3436) );
  CND3XL U2730 ( .A(n2719), .B(n3441), .C(n3440), .Z(n813) );
  CANR1XL U2731 ( .A(result[13]), .B(n2891), .C(n3439), .Z(n3440) );
  CND3XL U2732 ( .A(n2881), .B(n3517), .C(n3438), .Z(n3441) );
  CND3XL U2733 ( .A(n2743), .B(n3449), .C(n3448), .Z(n809) );
  CANR1XL U2734 ( .A(result[17]), .B(n2891), .C(n3447), .Z(n3448) );
  CND3XL U2735 ( .A(n2648), .B(n3490), .C(n3489), .Z(n824) );
  CANR1XL U2736 ( .A(result[2]), .B(n2891), .C(n3488), .Z(n3489) );
  CND3XL U2737 ( .A(n2662), .B(n3495), .C(n3494), .Z(n822) );
  CANR1XL U2738 ( .A(result[4]), .B(n2891), .C(n3493), .Z(n3494) );
  CND3XL U2739 ( .A(n2686), .B(n3504), .C(n3503), .Z(n818) );
  CANR1XL U2740 ( .A(result[8]), .B(n2891), .C(n3502), .Z(n3503) );
  CND3XL U2741 ( .A(n2700), .B(n3509), .C(n3508), .Z(n816) );
  CANR1XL U2742 ( .A(result[10]), .B(n2891), .C(n3507), .Z(n3508) );
  CND3XL U2743 ( .A(n2724), .B(n3521), .C(n3520), .Z(n812) );
  CANR1XL U2744 ( .A(result[14]), .B(n2891), .C(n3519), .Z(n3520) );
  CND3XL U2745 ( .A(n2738), .B(n3527), .C(n3526), .Z(n810) );
  CANR1XL U2746 ( .A(result[16]), .B(n2891), .C(n3525), .Z(n3526) );
  CND3XL U2747 ( .A(n2167), .B(n2166), .C(n2168), .Z(n953) );
  COR4X1 U2748 ( .A(n2154), .B(n3060), .C(i[5]), .D(n2171), .Z(n2167) );
  CND3XL U2749 ( .A(n2693), .B(n3433), .C(n3432), .Z(n817) );
  CANR1XL U2750 ( .A(result[9]), .B(n2891), .C(n3431), .Z(n3432) );
  CND3XL U2751 ( .A(n2881), .B(n3505), .C(n3430), .Z(n3433) );
  CND3XL U2752 ( .A(n2731), .B(n3445), .C(n3444), .Z(n811) );
  CANR1XL U2753 ( .A(result[15]), .B(n2891), .C(n3443), .Z(n3444) );
  CND3XL U2754 ( .A(n2881), .B(n3523), .C(n3442), .Z(n3445) );
  CND3XL U2755 ( .A(n2769), .B(n3458), .C(n3457), .Z(n805) );
  CANR1XL U2756 ( .A(result[21]), .B(n2891), .C(n3456), .Z(n3457) );
  CND3XL U2757 ( .A(n2881), .B(n3541), .C(n3455), .Z(n3458) );
  CND3XL U2758 ( .A(n2781), .B(n3462), .C(n3461), .Z(n803) );
  CANR1XL U2759 ( .A(result[23]), .B(n2891), .C(n3460), .Z(n3461) );
  CND3XL U2760 ( .A(n2795), .B(n3469), .C(n3468), .Z(n801) );
  CANR1XL U2761 ( .A(result[25]), .B(n2891), .C(n3467), .Z(n3468) );
  CND3XL U2762 ( .A(n2881), .B(n3554), .C(n3466), .Z(n3469) );
  CND3XL U2763 ( .A(n2807), .B(n3475), .C(n3474), .Z(n799) );
  CANR1XL U2764 ( .A(result[27]), .B(n2891), .C(n3473), .Z(n3474) );
  CND3XL U2765 ( .A(n2881), .B(n3559), .C(n3472), .Z(n3475) );
  CND3XL U2766 ( .A(n2819), .B(n3480), .C(n3479), .Z(n797) );
  CANR1XL U2767 ( .A(result[29]), .B(n2891), .C(n3478), .Z(n3479) );
  CND3XL U2768 ( .A(n2674), .B(n3499), .C(n3498), .Z(n820) );
  CANR1XL U2769 ( .A(result[6]), .B(n2891), .C(n3497), .Z(n3498) );
  CND3XL U2770 ( .A(n2712), .B(n3515), .C(n3514), .Z(n814) );
  CANR1XL U2771 ( .A(result[12]), .B(n2891), .C(n3513), .Z(n3514) );
  CND3XL U2772 ( .A(n2881), .B(n3512), .C(n3511), .Z(n3515) );
  CND3XL U2773 ( .A(n2750), .B(n3534), .C(n3533), .Z(n808) );
  CANR1XL U2774 ( .A(result[18]), .B(n2891), .C(n3532), .Z(n3533) );
  CND3XL U2775 ( .A(n2881), .B(n3531), .C(n3530), .Z(n3534) );
  CND3XL U2776 ( .A(n2762), .B(n3539), .C(n3538), .Z(n806) );
  CANR1XL U2777 ( .A(result[20]), .B(n2891), .C(n3537), .Z(n3538) );
  CND3XL U2778 ( .A(n2776), .B(n3545), .C(n3544), .Z(n804) );
  CANR1XL U2779 ( .A(result[22]), .B(n2891), .C(n3543), .Z(n3544) );
  CND3XL U2780 ( .A(n2788), .B(n3552), .C(n3551), .Z(n802) );
  CANR1XL U2781 ( .A(result[24]), .B(n2891), .C(n3550), .Z(n3551) );
  CND3XL U2782 ( .A(n2881), .B(n3549), .C(n3548), .Z(n3552) );
  CND3XL U2783 ( .A(n2800), .B(n3558), .C(n3557), .Z(n800) );
  CANR1XL U2784 ( .A(result[26]), .B(n2891), .C(n3556), .Z(n3557) );
  CND2X1 U2785 ( .A(n3051), .B(n2802), .Z(n2800) );
  CND3XL U2786 ( .A(n2814), .B(n3563), .C(n3562), .Z(n798) );
  CANR1XL U2787 ( .A(result[28]), .B(n2891), .C(n3561), .Z(n3562) );
  CND3XL U2788 ( .A(n2826), .B(n3570), .C(n3569), .Z(n796) );
  CANR1XL U2789 ( .A(result[30]), .B(n2891), .C(n3568), .Z(n3569) );
  CND3XL U2790 ( .A(n2881), .B(n3567), .C(n3566), .Z(n3570) );
  CAN2X1 U2791 ( .A(res_not_wire[44]), .B(n2901), .Z(n3013) );
  CENX1 U2792 ( .A(result[54]), .B(n3222), .Z(n3014) );
  COR2X1 U2793 ( .A(n3015), .B(n3700), .Z(n3392) );
  CND2IX1 U2794 ( .B(n3486), .A(n3072), .Z(n3417) );
  CND2IX1 U2795 ( .B(i[31]), .A(n2853), .Z(n2846) );
  CANR1XL U2796 ( .A(result[52]), .B(n3754), .C(n3670), .Z(n3671) );
  CNR2IX1 U2797 ( .B(result[18]), .A(n3046), .Z(n3451) );
  CNR2IX1 U2798 ( .B(result[30]), .A(n3047), .Z(n3483) );
  CND2X1 U2799 ( .A(res_not_wire[36]), .B(res_not_wire[32]), .Z(n3085) );
  CNR2X1 U2800 ( .A(n126), .B(n3058), .Z(n3363) );
  CNR2IX1 U2801 ( .B(n2901), .A(n3058), .Z(n3609) );
  CNR2IX1 U2802 ( .B(n3697), .A(n3058), .Z(n3699) );
  CANR2X1 U2803 ( .A(result[24]), .B(n3055), .C(n3053), .D(n2067), .Z(n2275)
         );
  CNR2IX1 U2804 ( .B(n3748), .A(n3058), .Z(n3724) );
  CNR2IX1 U2805 ( .B(res_not_wire[44]), .A(n3058), .Z(n3726) );
  CNR2IX1 U2806 ( .B(res_not_wire[40]), .A(n3058), .Z(n3354) );
  CANR2X1 U2807 ( .A(result[18]), .B(n3056), .C(n3054), .D(n2070), .Z(n2269)
         );
  CNR2IX1 U2808 ( .B(res_not_wire[6]), .A(n3058), .Z(n3356) );
  CANR2X1 U2809 ( .A(result[6]), .B(n3055), .C(n3052), .D(n2076), .Z(n2257) );
  CNR2IX1 U2810 ( .B(res_not_wire[38]), .A(n3058), .Z(n3358) );
  CNR2IX1 U2811 ( .B(res_not_wire[42]), .A(n3058), .Z(n3360) );
  CANR2X1 U2812 ( .A(result[12]), .B(n3056), .C(n3053), .D(n2073), .Z(n2263)
         );
  COND1XL U2813 ( .A(n3482), .B(n134), .C(n3370), .Z(n3371) );
  COND1XL U2814 ( .A(n3750), .B(n3577), .C(n130), .Z(n3578) );
  CND2X1 U2815 ( .A(n3662), .B(n3661), .Z(n838) );
  CANR1XL U2816 ( .A(result[51]), .B(n3754), .C(n3660), .Z(n3661) );
  CANR1XL U2817 ( .A(result[56]), .B(n3754), .C(n3694), .Z(n3695) );
  CND2X1 U2818 ( .A(n3583), .B(n3582), .Z(n853) );
  CANR1XL U2819 ( .A(result[36]), .B(n3754), .C(n3581), .Z(n3582) );
  CNR2X1 U2820 ( .A(n3580), .B(n2898), .Z(n3583) );
  CANR1XL U2821 ( .A(n3704), .B(n3587), .C(n3586), .Z(n3590) );
  CANR1XL U2822 ( .A(result[35]), .B(n3754), .C(n3588), .Z(n3589) );
  CND2X1 U2823 ( .A(n3598), .B(n3597), .Z(n842) );
  CANR1XL U2824 ( .A(result[47]), .B(n3754), .C(n3596), .Z(n3597) );
  CND2X1 U2825 ( .A(n3607), .B(n3606), .Z(n841) );
  CANR1XL U2826 ( .A(result[48]), .B(n3754), .C(n3605), .Z(n3606) );
  CNR2X1 U2827 ( .A(n3604), .B(n2987), .Z(n3607) );
  CND2X1 U2828 ( .A(n3617), .B(n3616), .Z(n851) );
  CANR1XL U2829 ( .A(result[38]), .B(n3754), .C(n3615), .Z(n3616) );
  CANR1XL U2830 ( .A(n3704), .B(n3628), .C(n3627), .Z(n3631) );
  CANR1XL U2831 ( .A(result[40]), .B(n3754), .C(n3629), .Z(n3630) );
  CND2X1 U2832 ( .A(n3643), .B(n3642), .Z(n847) );
  CANR1XL U2833 ( .A(result[42]), .B(n3754), .C(n3641), .Z(n3642) );
  CNR2X1 U2834 ( .A(n3640), .B(n2988), .Z(n3643) );
  CANR1XL U2835 ( .A(result[45]), .B(n3754), .C(n3650), .Z(n3651) );
  CND2X1 U2836 ( .A(n3685), .B(n3684), .Z(n835) );
  CANR1XL U2837 ( .A(result[54]), .B(n3754), .C(n3683), .Z(n3684) );
  CNR2X1 U2838 ( .A(n3682), .B(n2989), .Z(n3685) );
  CANR1XL U2839 ( .A(result[58]), .B(n3754), .C(n3717), .Z(n3718) );
  CANR1XL U2840 ( .A(n2881), .B(n3716), .C(n3715), .Z(n3719) );
  CANR1XL U2841 ( .A(result[39]), .B(n3754), .C(n3735), .Z(n3736) );
  CND2X1 U2842 ( .A(n3756), .B(n3755), .Z(n855) );
  CANR1XL U2843 ( .A(result[34]), .B(n3754), .C(n3753), .Z(n3755) );
  CNR2X1 U2844 ( .A(n3751), .B(n2990), .Z(n3756) );
  CND2X1 U2845 ( .A(n3351), .B(n3350), .Z(n834) );
  CANR1XL U2846 ( .A(result[55]), .B(n3754), .C(n3349), .Z(n3350) );
  CANR1XL U2847 ( .A(result[57]), .B(n3754), .C(n3251), .Z(n3252) );
  CANR1XL U2848 ( .A(result[37]), .B(n3754), .C(n3266), .Z(n3267) );
  CND2X1 U2849 ( .A(n3276), .B(n3275), .Z(n848) );
  CANR1XL U2850 ( .A(result[41]), .B(n3754), .C(n3274), .Z(n3275) );
  CENX1 U2851 ( .A(res_not_wire[40]), .B(n3043), .Z(n3272) );
  CANR1XL U2852 ( .A(result[43]), .B(n3754), .C(n3282), .Z(n3283) );
  CND2X1 U2853 ( .A(n3294), .B(n3293), .Z(n845) );
  CANR1XL U2854 ( .A(result[44]), .B(n3754), .C(n3292), .Z(n3293) );
  CANR1XL U2855 ( .A(n3704), .B(n3296), .C(n3295), .Z(n3299) );
  CANR1XL U2856 ( .A(result[46]), .B(n3754), .C(n3297), .Z(n3298) );
  CANR1XL U2857 ( .A(result[49]), .B(n3754), .C(n3307), .Z(n3308) );
  CNR2X1 U2858 ( .A(n3024), .B(n3306), .Z(n3309) );
  CANR1XL U2859 ( .A(result[50]), .B(n3754), .C(n3316), .Z(n3317) );
  CANR1XL U2860 ( .A(result[53]), .B(n3754), .C(n3332), .Z(n3333) );
  CANR2X1 U2861 ( .A(n3331), .B(n3330), .C(n2881), .D(n3329), .Z(n3334) );
  CND2X1 U2862 ( .A(n2179), .B(n2180), .Z(n947) );
  COR4X1 U2863 ( .A(n2153), .B(n3060), .C(i[7]), .D(n2176), .Z(n2180) );
  CND2X1 U2864 ( .A(n2184), .B(n2185), .Z(n945) );
  COND4CX1 U2865 ( .A(n2161), .B(n2011), .C(n2183), .D(i[9]), .Z(n2184) );
  CIVX2 U2866 ( .A(res_not_wire[14]), .Z(n3036) );
  CENX1 U2867 ( .A(opera1[24]), .B(n2900), .Z(n3186) );
  CND2X1 U2868 ( .A(i[14]), .B(n2198), .Z(n2197) );
  CND3XL U2869 ( .A(n1106), .B(n2102), .C(n56), .Z(n2235) );
  CEOX1 U2870 ( .A(result[48]), .B(n3207), .Z(n3599) );
  CEOXL U2871 ( .A(n3656), .B(n116), .Z(n3314) );
  CEOX1 U2872 ( .A(n3035), .B(res_not_wire[46]), .Z(n3594) );
  CENX1 U2873 ( .A(opera1[23]), .B(n2900), .Z(n3183) );
  CENX1 U2874 ( .A(opera1[22]), .B(n2900), .Z(n3191) );
  CNR3XL U2875 ( .A(n3764), .B(n56), .C(n2102), .Z(n2842) );
  CND2X1 U2876 ( .A(i[12]), .B(n2193), .Z(n2192) );
  CND2X1 U2877 ( .A(i[26]), .B(n2225), .Z(n2224) );
  COND11X1 U2878 ( .A(n2204), .B(i[18]), .C(n3060), .D(n2205), .Z(n936) );
  CND2X1 U2879 ( .A(i[18]), .B(n2206), .Z(n2205) );
  COND11X1 U2880 ( .A(n2209), .B(i[20]), .C(n3060), .D(n2210), .Z(n934) );
  COND2X1 U2881 ( .A(n1987), .B(n2147), .C(i[21]), .D(n2212), .Z(n933) );
  CENX1 U2882 ( .A(opera1[21]), .B(n2900), .Z(n3208) );
  CND3XL U2883 ( .A(i[19]), .B(i[18]), .C(n2007), .Z(n2209) );
  CND3XL U2884 ( .A(n3059), .B(i[20]), .C(n2005), .Z(n2212) );
  COR2X1 U2885 ( .A(n3026), .B(n3181), .Z(n3301) );
  CND3XL U2886 ( .A(n53), .B(n2170), .C(n56), .Z(n2166) );
  COND1XL U2887 ( .A(n2101), .B(n2908), .C(n2155), .Z(n957) );
  CANR2X1 U2888 ( .A(n3757), .B(n1998), .C(nst[0]), .D(n2157), .Z(n2155) );
  COND1XL U2889 ( .A(n2235), .B(n2004), .C(n2239), .Z(n921) );
  CANR2X1 U2890 ( .A(n3757), .B(n1998), .C(nst[2]), .D(n2157), .Z(n2239) );
  CND2X1 U2891 ( .A(n2199), .B(n2200), .Z(n939) );
  COR4X1 U2892 ( .A(n2150), .B(n3060), .C(i[15]), .D(n2196), .Z(n2200) );
  CND2X1 U2893 ( .A(n2221), .B(n2222), .Z(n929) );
  COR4X1 U2894 ( .A(n2092), .B(n3060), .C(i[25]), .D(n2218), .Z(n2222) );
  CND2X1 U2895 ( .A(n2226), .B(n2227), .Z(n927) );
  COND4CX1 U2896 ( .A(n3059), .B(n2095), .C(n2225), .D(i[27]), .Z(n2226) );
  CND2X1 U2897 ( .A(n2189), .B(n2190), .Z(n943) );
  COR4X1 U2898 ( .A(n2152), .B(n3060), .C(i[11]), .D(n2186), .Z(n2190) );
  CND2X1 U2899 ( .A(n2194), .B(n2195), .Z(n941) );
  CND2X1 U2900 ( .A(n2207), .B(n2208), .Z(n935) );
  CND2X1 U2901 ( .A(i[10]), .B(n2188), .Z(n2187) );
  CND2X1 U2902 ( .A(i[24]), .B(n2220), .Z(n2219) );
  CENX1 U2903 ( .A(n3505), .B(n3037), .Z(n3506) );
  CENX1 U2904 ( .A(opera1[25]), .B(n2900), .Z(n3108) );
  CENX1 U2905 ( .A(opera1[26]), .B(n2900), .Z(n3106) );
  CENX1 U2906 ( .A(opera1[27]), .B(n2900), .Z(n3103) );
  CENX1 U2907 ( .A(opera1[29]), .B(n2900), .Z(n3385) );
  COND1XL U2908 ( .A(n3517), .B(n152), .C(n3036), .Z(n3442) );
  COND1XL U2909 ( .A(n3554), .B(n140), .C(n3471), .Z(n3472) );
  COND1XL U2910 ( .A(n3547), .B(n3546), .C(n142), .Z(n3548) );
  COR2X1 U2911 ( .A(n3027), .B(n3549), .Z(n3554) );
  COND1XL U2912 ( .A(n1998), .B(n2047), .C(n2238), .Z(n922) );
  CND2X1 U2913 ( .A(n3261), .B(n3260), .Z(n3747) );
  CNR2IX1 U2914 ( .B(n3259), .A(n3463), .Z(n3260) );
  CNR3XL U2915 ( .A(n134), .B(n3255), .C(n3370), .Z(n3256) );
  CND2X1 U2916 ( .A(valid), .B(n3757), .Z(n2240) );
  CENX1 U2917 ( .A(n162), .B(n3491), .Z(n3492) );
  CENX1 U2918 ( .A(opera1[28]), .B(n2900), .Z(n3378) );
  COND1XL U2919 ( .A(n3510), .B(n2116), .C(n154), .Z(n3511) );
  COND1XL U2920 ( .A(n3529), .B(n3528), .C(n148), .Z(n3530) );
  CEOX1 U2921 ( .A(opera1[30]), .B(n2900), .Z(n3029) );
  CNR2X1 U2922 ( .A(n2927), .B(nst[0]), .Z(n55) );
  CANR1XL U2923 ( .A(n3743), .B(n3742), .C(n3741), .Z(n3744) );
  CND2X1 U2924 ( .A(n3743), .B(n3364), .Z(n3155) );
  CND2X1 U2925 ( .A(n3144), .B(n3122), .Z(n3145) );
  CANR2X1 U2926 ( .A(result[31]), .B(n3055), .C(n3053), .D(n2146), .Z(n2282)
         );
  CANR1XL U2927 ( .A(result[31]), .B(n2891), .C(n3483), .Z(n3484) );
  COND1XL U2928 ( .A(n134), .B(n3058), .C(n2282), .Z(n888) );
  CND3XL U2929 ( .A(n2833), .B(n3485), .C(n3484), .Z(n795) );
  CANR1XL U2930 ( .A(n2881), .B(n3080), .C(n3079), .Z(n3081) );
  COND4CX1 U2931 ( .A(n2161), .B(n2006), .C(n2206), .D(i[19]), .Z(n2207) );
  COND4CX1 U2932 ( .A(n2161), .B(n2092), .C(n2220), .D(i[25]), .Z(n2221) );
  CND2X1 U2933 ( .A(n2161), .B(n2093), .Z(n2230) );
  COND4CX1 U2934 ( .A(n2161), .B(n2147), .C(n2213), .D(i[22]), .Z(n2214) );
  COND4CX1 U2935 ( .A(n2161), .B(n2003), .C(n2202), .D(i[23]), .Z(n2216) );
  CANR1XL U2936 ( .A(n2243), .B(n3768), .C(n2244), .Z(n2241) );
  CANR2X1 U2937 ( .A(n3704), .B(n3315), .C(n2881), .D(n3314), .Z(n3318) );
  COND1XL U2938 ( .A(n2009), .B(n3060), .C(n2170), .Z(n2193) );
  CIVXL U2939 ( .A(n3420), .Z(n3034) );
  CND2IXL U2940 ( .B(n3012), .A(n3124), .Z(n3125) );
  COND1XL U2941 ( .A(n3346), .B(n3345), .C(n3344), .Z(n3688) );
  CENX1 U2942 ( .A(opera1[20]), .B(n2900), .Z(n3194) );
  CENX1 U2943 ( .A(opera1[19]), .B(n2900), .Z(n3198) );
  CND4XL U2944 ( .A(n3116), .B(n3115), .C(n2986), .D(n2971), .Z(n3167) );
  CND3XL U2945 ( .A(n3148), .B(n2985), .C(n2971), .Z(n3141) );
  CND2X1 U2946 ( .A(n3148), .B(n3144), .Z(n3149) );
  CNR2XL U2947 ( .A(n3121), .B(n3120), .Z(n3122) );
  COND1XL U2948 ( .A(n146), .B(n3058), .C(n2270), .Z(n900) );
  CND3XL U2949 ( .A(res_not_wire[20]), .B(n3535), .C(n2876), .Z(n3541) );
  CNR2IX2 U2950 ( .B(n3091), .A(n3090), .Z(n3092) );
  CND2XL U2951 ( .A(n2000), .B(n2093), .Z(n2229) );
  CNR2IX1 U2952 ( .B(n3636), .A(n3044), .Z(n3640) );
  CND4XL U2953 ( .A(i[28]), .B(n3059), .C(n2094), .D(n2000), .Z(n2231) );
  COND1XL U2954 ( .A(n2086), .B(n3060), .C(n2170), .Z(n2183) );
  COND11XL U2955 ( .A(n3060), .B(i[6]), .C(n2176), .D(n2177), .Z(n948) );
  CNR2IXL U2956 ( .B(result[51]), .A(n3045), .Z(n3670) );
  CNR2IXL U2957 ( .B(result[33]), .A(n3045), .Z(n3753) );
  CNR2IXL U2958 ( .B(result[57]), .A(n3045), .Z(n3717) );
  CNR2IXL U2959 ( .B(result[53]), .A(n3045), .Z(n3683) );
  CNR2IXL U2960 ( .B(result[50]), .A(n3045), .Z(n3660) );
  CNR2IXL U2961 ( .B(result[44]), .A(n3752), .Z(n3650) );
  COND1XL U2962 ( .A(i[0]), .B(n3060), .C(n2170), .Z(n2173) );
  COR3XL U2963 ( .A(i[0]), .B(i[11]), .C(n2852), .Z(n2851) );
  CND3XL U2964 ( .A(n3419), .B(n3418), .C(n2655), .Z(n823) );
  CND3XL U2965 ( .A(n3417), .B(n3416), .C(n2881), .Z(n3418) );
  CIVX2 U2966 ( .A(n2887), .Z(n3050) );
  CND3XL U2967 ( .A(n2757), .B(n3453), .C(n3452), .Z(n807) );
  CND3XL U2968 ( .A(n2881), .B(n3454), .C(n3450), .Z(n3453) );
  CANR1XL U2969 ( .A(result[19]), .B(n2891), .C(n3451), .Z(n3452) );
  CIVX2 U2970 ( .A(n2887), .Z(n3051) );
  CANR2X1 U2971 ( .A(n3704), .B(n3595), .C(n2881), .D(n3594), .Z(n3598) );
  CANR2X1 U2972 ( .A(n3704), .B(n3614), .C(n2881), .D(n3613), .Z(n3617) );
  CANR2X1 U2973 ( .A(n3704), .B(n3693), .C(n2881), .D(n3692), .Z(n3696) );
  COND11XL U2974 ( .A(n3060), .B(i[4]), .C(n2171), .D(n2175), .Z(n949) );
  COND11XL U2975 ( .A(n3060), .B(i[10]), .C(n2186), .D(n2187), .Z(n944) );
  CNR2IX1 U2976 ( .B(result[42]), .A(n3047), .Z(n3282) );
  CNR2IXL U2977 ( .B(result[40]), .A(n3045), .Z(n3274) );
  CNR2IX1 U2978 ( .B(result[56]), .A(n3045), .Z(n3251) );
  COND4CX1 U2979 ( .A(n3059), .B(n2149), .C(n2202), .D(i[17]), .Z(n2203) );
  COND4CXL U2980 ( .A(n2161), .B(n2150), .C(n2198), .D(i[15]), .Z(n2199) );
  COND4CX1 U2981 ( .A(n2161), .B(n2151), .C(n2193), .D(i[13]), .Z(n2194) );
  COND4CX1 U2982 ( .A(n2161), .B(n2152), .C(n2188), .D(i[11]), .Z(n2189) );
  COND4CX1 U2983 ( .A(n2162), .B(n2163), .C(n2148), .D(n2164), .Z(n954) );
  COND1XL U2984 ( .A(n3321), .B(n3319), .C(n3676), .Z(n3320) );
  COND11XL U2985 ( .A(n3060), .B(i[24]), .C(n2218), .D(n2219), .Z(n930) );
  CND2X1 U2986 ( .A(n2695), .B(n3051), .Z(n2693) );
  CND2X1 U2987 ( .A(n2752), .B(n3051), .Z(n2750) );
  CND2X1 U2988 ( .A(n2733), .B(n3051), .Z(n2731) );
  CND2X1 U2989 ( .A(n3051), .B(n2835), .Z(n2833) );
  CND2X1 U2990 ( .A(n3050), .B(n2650), .Z(n2648) );
  CND2X1 U2991 ( .A(n3050), .B(n2910), .Z(n2662) );
  CND2X1 U2992 ( .A(n3050), .B(n2669), .Z(n2667) );
  COND1XL U2993 ( .A(n2002), .B(n3060), .C(n2170), .Z(n2220) );
  CEOXL U2994 ( .A(n2670), .B(n2671), .Z(n2669) );
  CEOXL U2995 ( .A(n2689), .B(n2690), .Z(n2688) );
  CIVX2 U2996 ( .A(n3039), .Z(n3040) );
  CNR2XL U2997 ( .A(n3088), .B(n148), .Z(n3041) );
  CND3XL U2998 ( .A(i[17]), .B(i[16]), .C(n2215), .Z(n2204) );
  CND3XL U2999 ( .A(n3310), .B(n3323), .C(n3326), .Z(n3226) );
  CANR1XL U3000 ( .A(n3178), .B(n3179), .C(n3177), .Z(n3182) );
  CND2XL U3001 ( .A(n3216), .B(n3215), .Z(n3223) );
  CND2XL U3002 ( .A(n3216), .B(n3196), .Z(n3197) );
  COND1XL U3003 ( .A(n3038), .B(n3058), .C(n2260), .Z(n910) );
  COND1XL U3004 ( .A(n3486), .B(n164), .C(n3415), .Z(n3416) );
  COND1XL U3005 ( .A(n2162), .B(n2096), .C(n2174), .Z(n950) );
  CND2XL U3006 ( .A(result[63]), .B(n3049), .Z(n3572) );
  CND2XL U3007 ( .A(n2161), .B(n2096), .Z(n2163) );
  CND4XL U3008 ( .A(i[1]), .B(n3059), .C(n2096), .D(i[0]), .Z(n2174) );
  CND2X1 U3009 ( .A(n3051), .B(n2688), .Z(n2686) );
  CND2X1 U3010 ( .A(n3051), .B(n2707), .Z(n2705) );
  CND2X1 U3011 ( .A(n3051), .B(n2702), .Z(n2700) );
  CND2X1 U3012 ( .A(n3051), .B(n2721), .Z(n2719) );
  CND2X1 U3013 ( .A(n3051), .B(n2726), .Z(n2724) );
  CND2X1 U3014 ( .A(n3051), .B(n2740), .Z(n2738) );
  CND2X1 U3015 ( .A(n3051), .B(n2745), .Z(n2743) );
  CANR2XL U3016 ( .A(n2891), .B(result[1]), .C(n3049), .D(result[0]), .Z(n2642) );
  CND2IXL U3017 ( .B(n2882), .A(n3700), .Z(n3708) );
  CEOXL U3018 ( .A(n2760), .B(n2754), .Z(n2759) );
  CEOXL U3019 ( .A(n2651), .B(n2953), .Z(n2650) );
  CEOXL U3020 ( .A(n2765), .B(n2766), .Z(n2764) );
  CEOXL U3021 ( .A(c_inop2), .B(n2646), .Z(n2645) );
  CND3XL U3022 ( .A(n2881), .B(n3392), .C(n3376), .Z(n3391) );
  COND1XL U3023 ( .A(n3731), .B(n128), .C(n3730), .Z(n3732) );
  CND2X2 U3024 ( .A(n3092), .B(n3500), .Z(n3731) );
  COND11XL U3025 ( .A(n3060), .B(i[1]), .C(n2089), .D(n2172), .Z(n951) );
  COND2XL U3026 ( .A(n2089), .B(n2170), .C(i[0]), .D(n3060), .Z(n952) );
  COND3XL U3027 ( .A(n3246), .B(n2882), .C(n3245), .D(n3244), .Z(n830) );
  CNR2IXL U3028 ( .B(result[41]), .A(n3045), .Z(n3641) );
  CNR2IXL U3029 ( .B(result[39]), .A(n3045), .Z(n3629) );
  CNR2IXL U3030 ( .B(result[37]), .A(n3045), .Z(n3615) );
  CNR2IXL U3031 ( .B(result[47]), .A(n3045), .Z(n3605) );
  CNR2IXL U3032 ( .B(result[46]), .A(n3045), .Z(n3596) );
  CNR2IXL U3033 ( .B(result[34]), .A(n3047), .Z(n3588) );
  CNR2IXL U3034 ( .B(result[35]), .A(n3045), .Z(n3581) );
  CNR2IXL U3035 ( .B(result[29]), .A(n3045), .Z(n3568) );
  CNR2IXL U3036 ( .B(result[27]), .A(n3046), .Z(n3561) );
  CANR11XL U3037 ( .A(n2165), .B(n2148), .C(n3059), .D(n1990), .Z(n2164) );
  CANR1XL U3038 ( .A(res_not_wire[58]), .B(n3016), .C(n1073), .Z(n3709) );
  CND3XL U3039 ( .A(n2881), .B(n3496), .C(n2907), .Z(n3499) );
  CND2IXL U3040 ( .B(res_not_wire[6]), .A(n3496), .Z(n3425) );
  CNR3XL U3041 ( .A(n2885), .B(n1048), .C(n2235), .Z(n2246) );
  COND11XL U3042 ( .A(n3060), .B(i[14]), .C(n2196), .D(n2197), .Z(n940) );
  COND11XL U3043 ( .A(n3060), .B(i[30]), .C(n2233), .D(n2234), .Z(n924) );
  CND2IXL U3044 ( .B(n2099), .A(n3049), .Z(n3375) );
  COND4CXL U3045 ( .A(n2161), .B(n2233), .C(n1989), .D(i[30]), .Z(n2234) );
  CANR2XL U3046 ( .A(result[2]), .B(n3049), .C(result[3]), .D(n2891), .Z(n3419) );
  COND1XL U3047 ( .A(n2008), .B(n3060), .C(n2170), .Z(n2198) );
  CND2IXL U3048 ( .B(n2882), .A(n3571), .Z(n3413) );
  CANR1XL U3049 ( .A(n1081), .B(n3402), .C(res_not_wire[62]), .Z(n3414) );
  CND2IXL U3050 ( .B(res_not_wire[42]), .A(n3639), .Z(n3277) );
  CND3XL U3051 ( .A(n2881), .B(n3426), .C(n3425), .Z(n3429) );
  CANR1XL U3052 ( .A(n2903), .B(n3691), .C(res_not_wire[56]), .Z(n3250) );
  COND1XL U3053 ( .A(n3656), .B(n116), .C(n3655), .Z(n3657) );
  CND3XL U3054 ( .A(res_not_wire[8]), .B(n3500), .C(n3039), .Z(n3505) );
  CND2XL U3055 ( .A(n3500), .B(n3041), .Z(n3463) );
  CNR3XL U3056 ( .A(n3113), .B(n3112), .C(n3111), .Z(n3116) );
  CENX1 U3057 ( .A(opera1[15]), .B(opera1[31]), .Z(n3178) );
  CANR4CXL U3058 ( .A(n2747), .B(n2746), .C(n2753), .D(n2754), .Z(n2752) );
  CEOXL U3059 ( .A(n2741), .B(n2735), .Z(n2740) );
  CEOXL U3060 ( .A(n2817), .B(n2811), .Z(n2816) );
  CEOXL U3061 ( .A(n2822), .B(n2823), .Z(n2821) );
  CEOXL U3062 ( .A(n2746), .B(n2747), .Z(n2745) );
  CANR4CXL U3063 ( .A(n2728), .B(n2727), .C(n2734), .D(n2735), .Z(n2733) );
  CANR4CXL U3064 ( .A(n2804), .B(n2803), .C(n2810), .D(n2811), .Z(n2809) );
  COND1XL U3065 ( .A(n3040), .B(n3058), .C(n2258), .Z(n912) );
  CND2IXL U3066 ( .B(res_not_wire[54]), .A(n3681), .Z(n3335) );
  CND2IXL U3067 ( .B(res_not_wire[48]), .A(n3603), .Z(n3300) );
  CNR2IXL U3068 ( .B(res_not_wire[16]), .A(n3088), .Z(n3077) );
  CENX1 U3069 ( .A(n3571), .B(n2106), .Z(n3573) );
  CEOXL U3070 ( .A(n1983), .B(n2900), .Z(n3591) );
  COND3XL U3071 ( .A(n3654), .B(n3327), .C(n3326), .D(n3325), .Z(n3330) );
  CEOXL U3072 ( .A(n2722), .B(n2716), .Z(n2721) );
  CEOXL U3073 ( .A(n2703), .B(n2697), .Z(n2702) );
  CEOXL U3074 ( .A(n2779), .B(n2773), .Z(n2778) );
  CANR4CXL U3075 ( .A(n2709), .B(n2708), .C(n2715), .D(n2716), .Z(n2714) );
  CANR4CXL U3076 ( .A(n2690), .B(n2689), .C(n2696), .D(n2697), .Z(n2695) );
  CANR4CXL U3077 ( .A(n2766), .B(n2765), .C(n2772), .D(n2773), .Z(n2771) );
  CENX1 U3078 ( .A(result[63]), .B(n3409), .Z(n3410) );
  CND2XL U3079 ( .A(n3014), .B(n3225), .Z(n3346) );
  CND2XL U3080 ( .A(n3199), .B(n3197), .Z(n3203) );
  CEOXL U3081 ( .A(n2684), .B(n2678), .Z(n2683) );
  CEOXL U3082 ( .A(n2665), .B(n2659), .Z(n2664) );
  CEOXL U3083 ( .A(n2798), .B(n2792), .Z(n2797) );
  CANR4CXL U3084 ( .A(n2671), .B(n2670), .C(n2677), .D(n2678), .Z(n2676) );
  CANR4CXL U3085 ( .A(n2785), .B(n2784), .C(n2791), .D(n2792), .Z(n2790) );
  CANR4CXL U3086 ( .A(n2823), .B(n2822), .C(n2829), .D(n2830), .Z(n2828) );
  CANR4CXL U3087 ( .A(n2651), .B(n2953), .C(n2658), .D(n2659), .Z(n2657) );
  CANR2X1 U3088 ( .A(n2830), .B(n1984), .C(n1982), .D(n2877), .Z(n2841) );
  CIVX2 U3089 ( .A(n2161), .Z(n3060) );
  CIVX2 U3090 ( .A(n3067), .Z(n3757) );
  CIVX2 U3091 ( .A(n2933), .Z(n3758) );
  CIVX2 U3092 ( .A(n2235), .Z(n3768) );
  CIVX2 U3093 ( .A(i[30]), .Z(n3061) );
  CIVX2 U3094 ( .A(result[63]), .Z(n3769) );
  CIVX2 U3095 ( .A(n1026), .Z(n2106) );
  CIVX2 U3096 ( .A(n2236), .Z(n3065) );
  CIVX2 U3097 ( .A(result[62]), .Z(n3762) );
  CIVX2 U3098 ( .A(result[60]), .Z(n2083) );
  CIVX2 U3099 ( .A(res_not_wire[60]), .Z(n3761) );
  CIVX2 U3100 ( .A(result[56]), .Z(n2144) );
  CIVX2 U3101 ( .A(result[54]), .Z(n2135) );
  CIVX2 U3102 ( .A(res_not_wire[54]), .Z(n3765) );
  CIVX2 U3103 ( .A(result[52]), .Z(n2136) );
  CIVX2 U3104 ( .A(result[49]), .Z(n2137) );
  CIVX2 U3105 ( .A(result[48]), .Z(n2138) );
  CIVX2 U3106 ( .A(res_not_wire[48]), .Z(n3766) );
  CIVX2 U3107 ( .A(result[47]), .Z(n3759) );
  CIVX2 U3108 ( .A(res_not_wire[30]), .Z(n3767) );
  CIVX2 U3109 ( .A(result[0]), .Z(n3763) );
  CND2IX1 U3110 ( .B(n2887), .A(n2840), .Z(n3083) );
  CIVX2 U3111 ( .A(n3069), .Z(n3740) );
  CMXI2X1 U3112 ( .A0(n3071), .A1(n3070), .S(n2099), .Z(n3082) );
  CIVX2 U3113 ( .A(n160), .Z(n3073) );
  CIVX2 U3114 ( .A(res_not_wire[2]), .Z(n3415) );
  CIVX2 U3115 ( .A(n3496), .Z(n3074) );
  CIVX2 U3116 ( .A(n144), .Z(n3540) );
  CIVX2 U3117 ( .A(n138), .Z(n3078) );
  CIVX2 U3118 ( .A(res_not_wire[56]), .Z(n3084) );
  CIVX2 U3119 ( .A(n112), .Z(n3679) );
  CND2IX1 U3120 ( .B(n130), .A(res_not_wire[34]), .Z(n3253) );
  CIVX2 U3121 ( .A(n3731), .Z(n3093) );
  CIVX2 U3122 ( .A(n128), .Z(n3612) );
  CIVX2 U3123 ( .A(n3637), .Z(n3094) );
  CIVX2 U3124 ( .A(n3601), .Z(n3095) );
  CIVX2 U3125 ( .A(n3131), .Z(n3114) );
  CIVX2 U3126 ( .A(n3121), .Z(n3146) );
  CIVX2 U3127 ( .A(n3175), .Z(n3177) );
  CIVX2 U3128 ( .A(n3174), .Z(n3102) );
  CIVX2 U3129 ( .A(n3644), .Z(n3172) );
  CIVX2 U3130 ( .A(n3118), .Z(n3123) );
  CIVX2 U3131 ( .A(n3145), .Z(n3139) );
  CIVX2 U3132 ( .A(n3127), .Z(n3126) );
  CIVX2 U3133 ( .A(n3141), .Z(n3129) );
  CIVX2 U3134 ( .A(n3137), .Z(n3135) );
  CIVX2 U3135 ( .A(n3160), .Z(n3140) );
  CIVX2 U3136 ( .A(result[36]), .Z(n3158) );
  CIVX2 U3137 ( .A(n3149), .Z(n3147) );
  CIVX2 U3138 ( .A(n3176), .Z(n3180) );
  CENX1 U3139 ( .A(n3181), .B(n3026), .Z(n3302) );
  CIVX2 U3140 ( .A(n3204), .Z(n3664) );
  CND2IX1 U3141 ( .B(result[53]), .A(n3211), .Z(n3212) );
  CIVX2 U3142 ( .A(n3220), .Z(n3690) );
  CIVX2 U3143 ( .A(n3224), .Z(n3324) );
  CIVX2 U3144 ( .A(n3254), .Z(n3257) );
  CAN2X1 U3145 ( .A(n3257), .B(n3256), .Z(n3261) );
  CND2IX1 U3146 ( .B(res_not_wire[36]), .A(n3579), .Z(n3262) );
  CIVX2 U3147 ( .A(n3593), .Z(n3305) );
  COND1X2 U3148 ( .A(n3305), .B(n3592), .C(n3304), .Z(n3341) );
  CIVX2 U3149 ( .A(n3341), .Z(n3600) );
  CND2IX1 U3150 ( .B(n3312), .A(n3311), .Z(n3673) );
  CENX1 U3151 ( .A(n3313), .B(n3322), .Z(n3315) );
  CND2IX1 U3152 ( .B(n3322), .A(n3321), .Z(n3654) );
  CIVX2 U3153 ( .A(n3337), .Z(n3689) );
  CIVX2 U3154 ( .A(n3338), .Z(n3340) );
  CIVX2 U3155 ( .A(n3688), .Z(n3347) );
  CIVX2 U3156 ( .A(res_not_wire[0]), .Z(n3352) );
  CMXI2X1 U3157 ( .A0(n3053), .A1(n3055), .S(result[40]), .Z(n3353) );
  CND2IX1 U3158 ( .B(n3354), .A(n3353), .Z(n879) );
  CND2IX1 U3159 ( .B(n3355), .A(n2269), .Z(n901) );
  CND2IX1 U3160 ( .B(n3356), .A(n2257), .Z(n913) );
  CMXI2X1 U3161 ( .A0(n3052), .A1(n3056), .S(result[38]), .Z(n3357) );
  CND2IX1 U3162 ( .B(n3358), .A(n3357), .Z(n881) );
  CMXI2X1 U3163 ( .A0(n3054), .A1(n3057), .S(result[42]), .Z(n3359) );
  CND2IX1 U3164 ( .B(n3360), .A(n3359), .Z(n877) );
  CND2IX1 U3165 ( .B(n3361), .A(n2263), .Z(n907) );
  CMXI2X1 U3166 ( .A0(n3053), .A1(n3055), .S(result[39]), .Z(n3362) );
  CND2IX1 U3167 ( .B(n3363), .A(n3362), .Z(n880) );
  CIVX2 U3168 ( .A(n3365), .Z(n3741) );
  CMXI2X1 U3169 ( .A0(n3368), .A1(n3367), .S(n3366), .Z(n3374) );
  CIVX2 U3170 ( .A(n3701), .Z(n3384) );
  CENX1 U3171 ( .A(n1081), .B(n3402), .Z(n3400) );
  CENX1 U3172 ( .A(result[62]), .B(n3029), .Z(n3393) );
  COND3X1 U3173 ( .A(n3400), .B(n2882), .C(n3399), .D(n3398), .Z(n827) );
  CAN2X1 U3174 ( .A(res_not_wire[62]), .B(n1081), .Z(n3401) );
  CIVX2 U3175 ( .A(n3404), .Z(n3405) );
  CENX1 U3176 ( .A(res_not_wire[16]), .B(n3529), .Z(n3446) );
  CIVX2 U3177 ( .A(n3454), .Z(n3535) );
  CENX1 U3178 ( .A(res_not_wire[22]), .B(n3547), .Z(n3459) );
  CIVX2 U3179 ( .A(res_not_wire[26]), .Z(n3471) );
  CND2IX1 U3180 ( .B(res_not_wire[30]), .A(n3567), .Z(n3481) );
  CENX1 U3181 ( .A(n3517), .B(n3516), .Z(n3518) );
  CENX1 U3182 ( .A(n3523), .B(n3522), .Z(n3524) );
  CIVX2 U3183 ( .A(res_not_wire[16]), .Z(n3528) );
  CIVX2 U3184 ( .A(res_not_wire[22]), .Z(n3546) );
  CENX1 U3185 ( .A(n3554), .B(n3553), .Z(n3555) );
  CIVX2 U3186 ( .A(n3574), .Z(n3576) );
  CIVX2 U3187 ( .A(res_not_wire[34]), .Z(n3577) );
  CMXI2X1 U3188 ( .A0(n3052), .A1(n3056), .S(result[43]), .Z(n3608) );
  CND2IX1 U3189 ( .B(n3609), .A(n3608), .Z(n876) );
  CIVX2 U3190 ( .A(n3621), .Z(n3622) );
  CMXI2X1 U3191 ( .A0(n3626), .A1(n3625), .S(n3011), .Z(n3628) );
  CIVX2 U3192 ( .A(res_not_wire[50]), .Z(n3655) );
  CIVX2 U3193 ( .A(n3663), .Z(n3666) );
  CIVX2 U3194 ( .A(n3686), .Z(n3687) );
  CMXI2X1 U3195 ( .A0(n3054), .A1(n3057), .S(result[45]), .Z(n3698) );
  CND2IX1 U3196 ( .B(n3699), .A(n3698), .Z(n874) );
  COND3X1 U3197 ( .A(n3709), .B(n3708), .C(n3707), .D(n3706), .Z(n829) );
  CND2IX1 U3198 ( .B(n3721), .A(n3720), .Z(n883) );
  CND2IX1 U3199 ( .B(n3722), .A(n2275), .Z(n895) );
  CND2IX1 U3200 ( .B(n3724), .A(n3723), .Z(n886) );
  CMXI2X1 U3201 ( .A0(n3053), .A1(n3056), .S(result[44]), .Z(n3725) );
  CND2IX1 U3202 ( .B(n3726), .A(n3725), .Z(n875) );
  CIVX2 U3203 ( .A(n3727), .Z(n3728) );
  CIVX2 U3204 ( .A(res_not_wire[38]), .Z(n3730) );
  CENX1 U3205 ( .A(n3739), .B(n3760), .Z(n3745) );
endmodule



module multiplier ( result, valid, opera1, opera2, muordi, clock, reset, start
 );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input muordi, clock, reset, start;
  output valid;
  wire   opera2_63, N34, n52, n53, n55, n56, n106, n110, n112, n114, n116,
         n118, n120, n122, n124, n126, n128, n130, n132, n134, n136, n138,
         n140, n142, n144, n146, n148, n150, n154, n158, n160, n162, n164,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n960, n962, n1053, n1056, n1061, n1093, n1119, n2001, n2002, n2003,
         n2004, n2005, n2007, n2008, n2015, n2016, n2023, n2029, n2031, n2032,
         n2033, n2034, n2035, n2036, n2038, n2040, n2042, n2044, n2045, n2046,
         n2047, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2085, n2086, n2088, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2110, n2112, n2113, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2129, n2130,
         n2133, n2137, n2138, n2140, n2141, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2159, n2162, n2163, n2164, n2166, n2167, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2297, n2298, n2300,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2330, n2347, n2348, n2630, n2631, n2633,
         n2634, n2635, n2637, n2638, n2639, n2642, n2643, n2644, n2645, n2646,
         n2649, n2650, n2651, n2652, n2653, n2655, n2656, n2657, n2658, n2661,
         n2662, n2663, n2664, n2665, n2668, n2669, n2670, n2671, n2672, n2674,
         n2675, n2676, n2677, n2680, n2681, n2682, n2683, n2684, n2687, n2688,
         n2689, n2690, n2691, n2693, n2694, n2695, n2696, n2699, n2700, n2701,
         n2702, n2703, n2706, n2707, n2708, n2709, n2710, n2712, n2713, n2714,
         n2715, n2718, n2719, n2720, n2721, n2722, n2725, n2726, n2727, n2728,
         n2729, n2731, n2732, n2733, n2734, n2737, n2738, n2739, n2740, n2741,
         n2744, n2745, n2746, n2747, n2748, n2750, n2751, n2752, n2753, n2756,
         n2757, n2758, n2759, n2760, n2763, n2764, n2766, n2767, n2769, n2770,
         n2771, n2772, n2775, n2776, n2777, n2778, n2779, n2782, n2783, n2785,
         n2786, n2788, n2789, n2790, n2791, n2794, n2795, n2796, n2797, n2798,
         n2801, n2802, n2803, n2804, n2805, n2807, n2808, n2809, n2810, n2813,
         n2814, n2815, n2816, n2817, n2820, n2821, n2823, n2824, n2826, n2829,
         n2833, n2834, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703;
  wire   [63:0] res_not_wire;
  wire   [2:0] nst;
  wire   [31:0] i;
  tri   c_inop1;
  tri   c_inop2;
  tri   c_inres;
  assign opera2_63 = opera2[63];

  CTSX2 A4 ( .A(1'b0), .E(n2002), .Z(c_inop2) );
  CTSX2 A3 ( .A(1'b1), .E(opera2_63), .Z(c_inop2) );
  CTSX2 A6 ( .A(1'b0), .E(n2137), .Z(c_inres) );
  CTSX2 A5 ( .A(1'b1), .E(n1061), .Z(c_inres) );
  CIVX2 U1667 ( .A(n2821), .Z(n2001) );
  CIVX2 U1670 ( .A(n2167), .Z(n2004) );
  CIVX2 U1671 ( .A(n2204), .Z(n2005) );
  CIVX2 U1673 ( .A(n2178), .Z(n2007) );
  CIVX2 U1674 ( .A(n2174), .Z(n2008) );
  CIVX2 U1681 ( .A(reset), .Z(n2015) );
  CIVX2 U1682 ( .A(n2166), .Z(n2016) );
  CIVX2 U1697 ( .A(res_not_wire[62]), .Z(n2031) );
  CIVX2 U1708 ( .A(result[37]), .Z(n2042) );
  CIVX2 U1711 ( .A(result[41]), .Z(n2045) );
  CIVX2 U1717 ( .A(result[31]), .Z(n2051) );
  CIVX2 U1719 ( .A(result[29]), .Z(n2053) );
  CIVX2 U1734 ( .A(result[30]), .Z(n2068) );
  CIVX2 U1754 ( .A(res_not_wire[48]), .Z(n2088) );
  CIVX2 U1756 ( .A(res_not_wire[54]), .Z(n2090) );
  CIVX2 U1761 ( .A(res_not_wire[42]), .Z(n2095) );
  CIVX2 U1767 ( .A(n2255), .Z(n2101) );
  CIVX2 U1771 ( .A(n2227), .Z(n2105) );
  CIVX2 U1783 ( .A(n2222), .Z(n2117) );
  CIVX2 U1784 ( .A(n2217), .Z(n2118) );
  CIVX2 U1790 ( .A(res_not_wire[24]), .Z(n2124) );
  CIVX2 U1791 ( .A(res_not_wire[18]), .Z(n2125) );
  CIVX2 U1796 ( .A(n2212), .Z(n2130) );
  CIVX2 U1804 ( .A(res_not_wire[0]), .Z(n2138) );
  CIVX2 U1806 ( .A(n2834), .Z(n2140) );
  CIVX2 U1807 ( .A(n53), .Z(n2141) );
  CIVX2 U1809 ( .A(i[8]), .Z(n2143) );
  CIVX2 U1810 ( .A(n2207), .Z(n2144) );
  CIVX2 U1812 ( .A(n2195), .Z(n2146) );
  CIVX2 U1814 ( .A(n2190), .Z(n2148) );
  CIVX2 U1815 ( .A(n2185), .Z(n2149) );
  CIVX2 U1818 ( .A(n2180), .Z(n2150) );
  CIVX2 U1827 ( .A(n962), .Z(n2159) );
  CAOR2X1 U1832 ( .A(i[31]), .B(n2007), .C(n2169), .D(n3044), .Z(n955) );
  COR4X1 U1833 ( .A(n2155), .B(n3043), .C(i[5]), .D(n2180), .Z(n2175) );
  COR4X1 U1834 ( .A(n2163), .B(n3043), .C(i[7]), .D(n2185), .Z(n2189) );
  COR4X1 U1835 ( .A(n2143), .B(n3043), .C(i[9]), .D(n2190), .Z(n2194) );
  COR4X1 U1836 ( .A(n2154), .B(n3043), .C(i[11]), .D(n2195), .Z(n2199) );
  CND2IX1 U1837 ( .B(n2202), .A(i[12]), .Z(n2201) );
  COR4X1 U1838 ( .A(n2153), .B(n3043), .C(i[13]), .D(n2200), .Z(n2203) );
  COR4X1 U1839 ( .A(n2129), .B(n3043), .C(i[16]), .D(n2207), .Z(n2211) );
  COR4X1 U1840 ( .A(n2119), .B(n3043), .C(i[18]), .D(n2212), .Z(n2216) );
  COR4X1 U1841 ( .A(n2123), .B(n3043), .C(i[20]), .D(n2217), .Z(n2221) );
  COR4X1 U1842 ( .A(n2122), .B(n3043), .C(i[22]), .D(n2222), .Z(n2226) );
  COR2X1 U1843 ( .A(i[24]), .B(n2227), .Z(n2230) );
  CND2IX1 U1844 ( .B(n2234), .A(n2103), .Z(n2233) );
  COR4X1 U1845 ( .A(n2103), .B(n3043), .C(i[26]), .D(n2234), .Z(n2236) );
  COR4X1 U1846 ( .A(n3043), .B(n2102), .C(n2100), .D(i[28]), .Z(n2240) );
  CAOR2X1 U1847 ( .A(valid), .B(n2857), .C(n3034), .D(n3701), .Z(n923) );
  CAN4X1 U1848 ( .A(n2249), .B(n2252), .C(n2253), .D(n2254), .Z(n2166) );
  CAN4X1 U1874 ( .A(n56), .B(n53), .C(n1119), .D(reset), .Z(n2256) );
  CNR8X1 U1875 ( .A(i[1]), .B(i[19]), .C(i[16]), .D(i[2]), .E(n2839), .F(n2840), .G(n2837), .H(n2841), .Z(n2255) );
  COR3X1 U1876 ( .A(i[0]), .B(i[11]), .C(n2842), .Z(n2841) );
  COR6X1 U1877 ( .A(i[11]), .B(n2842), .C(n2840), .D(i[5]), .E(i[19]), .F(
        i[16]), .Z(n2843) );
  COR8X1 U1878 ( .A(i[20]), .B(i[17]), .C(i[22]), .D(i[21]), .E(i[26]), .F(
        i[24]), .G(i[9]), .H(i[30]), .Z(n2842) );
  COR8X1 U1879 ( .A(i[13]), .B(i[12]), .C(i[10]), .D(n2844), .E(i[28]), .F(
        i[27]), .G(i[25]), .H(n2845), .Z(n2840) );
  COR4X1 U1880 ( .A(i[29]), .B(i[6]), .C(i[7]), .D(i[8]), .Z(n2845) );
  COR4X1 U1881 ( .A(i[14]), .B(i[15]), .C(i[18]), .D(i[23]), .Z(n2844) );
  CND2IX1 U1882 ( .B(n2878), .A(nst[1]), .Z(n52) );
  CFD1XL \res_not_reg[54]  ( .D(n865), .CP(clock), .Q(res_not_wire[54]), .QN(
        n2959) );
  CFD1XL \res_not_reg[30]  ( .D(n889), .CP(clock), .Q(res_not_wire[30]), .QN(
        n2993) );
  CFD1QXL \result_reg[31]  ( .D(n794), .CP(clock), .Q(result[31]) );
  CFD1XL \res_not_reg[59]  ( .D(n860), .CP(clock), .QN(n106) );
  CFD1QXL \result_reg[29]  ( .D(n2876), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[30]  ( .D(n2877), .CP(clock), .Q(result[30]) );
  CFD1XL \res_not_reg[55]  ( .D(n864), .CP(clock), .QN(n110) );
  CFD1XL \res_not_reg[51]  ( .D(n868), .CP(clock), .QN(n114) );
  CFD1XL \res_not_reg[53]  ( .D(n866), .CP(clock), .Q(n2871), .QN(n112) );
  CFD1XL \res_not_reg[49]  ( .D(n870), .CP(clock), .QN(n116) );
  CFD1XL \res_not_reg[33]  ( .D(n886), .CP(clock), .Q(n2965), .QN(n132) );
  CFD1XL \res_not_reg[47]  ( .D(n872), .CP(clock), .QN(n118) );
  CFD1XL \res_not_reg[35]  ( .D(n884), .CP(clock), .QN(n130) );
  CFD1XL \res_not_reg[41]  ( .D(n878), .CP(clock), .QN(n124) );
  CFD1XL \res_not_reg[31]  ( .D(n888), .CP(clock), .Q(n2869), .QN(n134) );
  CFD1XL \res_not_reg[36]  ( .D(n883), .CP(clock), .Q(res_not_wire[36]), .QN(
        n2953) );
  CFD1XL \res_not_reg[37]  ( .D(n882), .CP(clock), .QN(n128) );
  CFD1XL \res_not_reg[43]  ( .D(n876), .CP(clock), .QN(n122) );
  CFD1XL \res_not_reg[23]  ( .D(n896), .CP(clock), .QN(n142) );
  CFD1XL \res_not_reg[25]  ( .D(n894), .CP(clock), .QN(n140) );
  CFD1XL \res_not_reg[29]  ( .D(n890), .CP(clock), .QN(n136) );
  CFD1XL \res_not_reg[27]  ( .D(n892), .CP(clock), .QN(n138) );
  CFD1XL \res_not_reg[45]  ( .D(n874), .CP(clock), .Q(n2870), .QN(n120) );
  CFD1XL \result_reg[49]  ( .D(n839), .CP(clock), .Q(result[49]), .QN(n2961)
         );
  CFD1XL \res_not_reg[21]  ( .D(n898), .CP(clock), .QN(n144) );
  CFD1XL \res_not_reg[17]  ( .D(n902), .CP(clock), .QN(n148) );
  CFD1XL \res_not_reg[19]  ( .D(n900), .CP(clock), .Q(n2868), .QN(n146) );
  CFD1XL \result_reg[48]  ( .D(n840), .CP(clock), .Q(result[48]), .QN(n2962)
         );
  CFD1XL \res_not_reg[11]  ( .D(n908), .CP(clock), .QN(n154) );
  CFD1XL \res_not_reg[15]  ( .D(n904), .CP(clock), .Q(n2867), .QN(n150) );
  CFD1XL \result_reg[38]  ( .D(n850), .CP(clock), .Q(result[38]), .QN(n2960)
         );
  CFD1XL \result_reg[39]  ( .D(n849), .CP(clock), .Q(result[39]), .QN(n2963)
         );
  CFD1XL \result_reg[40]  ( .D(n848), .CP(clock), .Q(result[40]), .QN(n2955)
         );
  CFD1XL \res_not_reg[4]  ( .D(n915), .CP(clock), .Q(res_not_wire[4]), .QN(
        n3002) );
  CFD1XL \res_not_reg[5]  ( .D(n914), .CP(clock), .QN(n160) );
  CFD1XL \res_not_reg[7]  ( .D(n912), .CP(clock), .Q(n2863), .QN(n158) );
  CTSX2 A2 ( .A(1'b0), .E(n2859), .Z(c_inop1) );
  CTSX2 A1 ( .A(1'b1), .E(opera1[31]), .Z(c_inop1) );
  CFD1XL \result_reg[35]  ( .D(n853), .CP(clock), .Q(result[35]), .QN(n2950)
         );
  CFD1QX1 \result_reg[61]  ( .D(n827), .CP(clock), .Q(result[61]) );
  CFD1XL \res_not_reg[3]  ( .D(n916), .CP(clock), .QN(n162) );
  CFD1XL \res_not_reg[0]  ( .D(n920), .CP(clock), .Q(res_not_wire[0]), .QN(
        n2932) );
  CFD1QXL \result_reg[63]  ( .D(n919), .CP(clock), .Q(result[63]) );
  CFD4QXL \cst_reg[0]  ( .D(n55), .CP(clock), .SD(n2015), .Q(n56) );
  CFD4QXL \cst_reg[1]  ( .D(n52), .CP(clock), .SD(n2015), .Q(n53) );
  CFD2XL \cst_reg[2]  ( .D(N34), .CP(clock), .CD(n2015), .Q(n3699), .QN(n1119)
         );
  CFD1XL \res_not_reg[39]  ( .D(n880), .CP(clock), .Q(n3226), .QN(n126) );
  CFD1X1 sign_reg ( .D(n2879), .CP(clock), .Q(n1061), .QN(n2137) );
  CFD1QXL valid_reg ( .D(n923), .CP(clock), .Q(valid) );
  CFD1QXL \i_reg[8]  ( .D(n946), .CP(clock), .Q(i[8]) );
  CFD1QXL \res_not_reg[38]  ( .D(n881), .CP(clock), .Q(res_not_wire[38]) );
  CFD1QXL \res_not_reg[32]  ( .D(n887), .CP(clock), .Q(res_not_wire[32]) );
  CFD1QXL \res_not_reg[2]  ( .D(n917), .CP(clock), .Q(res_not_wire[2]) );
  CFD1QXL \res_not_reg[14]  ( .D(n905), .CP(clock), .Q(res_not_wire[14]) );
  CFD1QXL \res_not_reg[13]  ( .D(n906), .CP(clock), .Q(n960) );
  CFD1QXL \res_not_reg[10]  ( .D(n909), .CP(clock), .Q(res_not_wire[10]) );
  CFD1QXL \res_not_reg[8]  ( .D(n911), .CP(clock), .Q(res_not_wire[8]) );
  CFD1QXL \res_not_reg[28]  ( .D(n891), .CP(clock), .Q(res_not_wire[28]) );
  CFD1QXL \res_not_reg[26]  ( .D(n893), .CP(clock), .Q(res_not_wire[26]) );
  CFD1QXL \res_not_reg[24]  ( .D(n895), .CP(clock), .Q(res_not_wire[24]) );
  CFD1QXL \res_not_reg[63]  ( .D(n793), .CP(clock), .Q(n1056) );
  CFD1QXL \res_not_reg[62]  ( .D(n857), .CP(clock), .Q(res_not_wire[62]) );
  CFD1QXL \res_not_reg[61]  ( .D(n858), .CP(clock), .Q(n1053) );
  CFD1QXL \res_not_reg[60]  ( .D(n859), .CP(clock), .Q(res_not_wire[60]) );
  CFD1QXL \res_not_reg[58]  ( .D(n861), .CP(clock), .Q(res_not_wire[58]) );
  CFD1QXL \res_not_reg[57]  ( .D(n862), .CP(clock), .Q(n1093) );
  CFD1QXL \res_not_reg[56]  ( .D(n863), .CP(clock), .Q(res_not_wire[56]) );
  CFD1QXL \res_not_reg[52]  ( .D(n867), .CP(clock), .Q(res_not_wire[52]) );
  CFD1QXL \res_not_reg[50]  ( .D(n869), .CP(clock), .Q(res_not_wire[50]) );
  CFD1QXL \res_not_reg[48]  ( .D(n871), .CP(clock), .Q(res_not_wire[48]) );
  CFD1QXL \res_not_reg[46]  ( .D(n873), .CP(clock), .Q(res_not_wire[46]) );
  CFD1QXL \res_not_reg[44]  ( .D(n875), .CP(clock), .Q(res_not_wire[44]) );
  CFD1QXL \res_not_reg[42]  ( .D(n877), .CP(clock), .Q(res_not_wire[42]) );
  CFD1QXL \res_not_reg[40]  ( .D(n879), .CP(clock), .Q(res_not_wire[40]) );
  CFD1QXL \res_not_reg[22]  ( .D(n897), .CP(clock), .Q(res_not_wire[22]) );
  CFD1QXL \res_not_reg[20]  ( .D(n899), .CP(clock), .Q(res_not_wire[20]) );
  CFD1QXL \res_not_reg[18]  ( .D(n901), .CP(clock), .Q(res_not_wire[18]) );
  CFD1QXL \res_not_reg[16]  ( .D(n903), .CP(clock), .Q(res_not_wire[16]) );
  CFD1QXL \res_not_reg[9]  ( .D(n910), .CP(clock), .Q(n962) );
  CFD1QXL \res_not_reg[6]  ( .D(n913), .CP(clock), .Q(res_not_wire[6]) );
  CFD1QXL \res_not_reg[34]  ( .D(n885), .CP(clock), .Q(res_not_wire[34]) );
  CFD1QXL \result_reg[47]  ( .D(n841), .CP(clock), .Q(result[47]) );
  CFD1QXL \result_reg[34]  ( .D(n854), .CP(clock), .Q(result[34]) );
  CFD1QXL \result_reg[36]  ( .D(n852), .CP(clock), .Q(result[36]) );
  CFD1QXL \result_reg[41]  ( .D(n847), .CP(clock), .Q(result[41]) );
  CFD1QXL \result_reg[52]  ( .D(n836), .CP(clock), .Q(result[52]) );
  CFD1QXL \result_reg[46]  ( .D(n842), .CP(clock), .Q(result[46]) );
  CFD1QXL \result_reg[37]  ( .D(n851), .CP(clock), .Q(result[37]) );
  CFD1QXL \result_reg[50]  ( .D(n838), .CP(clock), .Q(result[50]) );
  CFD1QXL \result_reg[42]  ( .D(n846), .CP(clock), .Q(result[42]) );
  CFD1QXL \result_reg[43]  ( .D(n845), .CP(clock), .Q(result[43]) );
  CFD1QXL \result_reg[51]  ( .D(n837), .CP(clock), .Q(result[51]) );
  CFD1QXL \result_reg[53]  ( .D(n835), .CP(clock), .Q(result[53]) );
  CFD1QXL \result_reg[54]  ( .D(n834), .CP(clock), .Q(result[54]) );
  CFD1QXL \result_reg[44]  ( .D(n844), .CP(clock), .Q(result[44]) );
  CFD1QXL \result_reg[57]  ( .D(n831), .CP(clock), .Q(result[57]) );
  CFD1QXL \result_reg[45]  ( .D(n843), .CP(clock), .Q(result[45]) );
  CFD1QXL \result_reg[55]  ( .D(n833), .CP(clock), .Q(result[55]) );
  CFD1QXL \result_reg[56]  ( .D(n832), .CP(clock), .Q(result[56]) );
  CFD1QXL \result_reg[59]  ( .D(n829), .CP(clock), .Q(result[59]) );
  CFD1QXL \result_reg[58]  ( .D(n830), .CP(clock), .Q(result[58]) );
  CFD1QXL \result_reg[60]  ( .D(n828), .CP(clock), .Q(result[60]) );
  CFD1XL \nst_reg[1]  ( .D(n2882), .CP(clock), .Q(nst[1]), .QN(n2049) );
  CFD1XL \nst_reg[2]  ( .D(n921), .CP(clock), .Q(nst[2]) );
  CFD1XL \nst_reg[0]  ( .D(n2884), .CP(clock), .Q(nst[0]) );
  CFD1XL \i_reg[0]  ( .D(n952), .CP(clock), .Q(i[0]), .QN(n2162) );
  CFD1XL \i_reg[1]  ( .D(n951), .CP(clock), .Q(i[1]), .QN(n2157) );
  CFD1XL \i_reg[23]  ( .D(n931), .CP(clock), .Q(i[23]), .QN(n2106) );
  CFD1XL \i_reg[21]  ( .D(n933), .CP(clock), .Q(i[21]), .QN(n2122) );
  CFD1XL \i_reg[19]  ( .D(n935), .CP(clock), .Q(i[19]), .QN(n2123) );
  CFD1XL \i_reg[17]  ( .D(n937), .CP(clock), .Q(i[17]), .QN(n2119) );
  CFD1XL \i_reg[15]  ( .D(n939), .CP(clock), .Q(i[15]), .QN(n2129) );
  CFD1XL \i_reg[10]  ( .D(n944), .CP(clock), .Q(i[10]), .QN(n2154) );
  CFD1XL \i_reg[4]  ( .D(n949), .CP(clock), .Q(i[4]), .QN(n2155) );
  CFD1XL \i_reg[25]  ( .D(n929), .CP(clock), .Q(i[25]), .QN(n2103) );
  CFD1XL \i_reg[22]  ( .D(n932), .CP(clock), .Q(i[22]) );
  CFD1XL \i_reg[7]  ( .D(n947), .CP(clock), .Q(i[7]) );
  CFD1XL \i_reg[6]  ( .D(n948), .CP(clock), .Q(i[6]), .QN(n2163) );
  CFD1XL \i_reg[27]  ( .D(n927), .CP(clock), .Q(i[27]), .QN(n2102) );
  CFD1XL \i_reg[20]  ( .D(n934), .CP(clock), .Q(i[20]) );
  CFD1XL \i_reg[18]  ( .D(n936), .CP(clock), .Q(i[18]) );
  CFD1XL \i_reg[9]  ( .D(n945), .CP(clock), .Q(i[9]) );
  CFD1XL \i_reg[5]  ( .D(n953), .CP(clock), .Q(i[5]) );
  CFD1XL \i_reg[16]  ( .D(n938), .CP(clock), .Q(i[16]) );
  CFD1XL \i_reg[11]  ( .D(n943), .CP(clock), .Q(i[11]) );
  CFD1XL \i_reg[26]  ( .D(n2886), .CP(clock), .Q(i[26]), .QN(n2121) );
  CFD1XL \i_reg[3]  ( .D(n954), .CP(clock), .Q(i[3]), .QN(n2151) );
  CFD1XL \i_reg[24]  ( .D(n930), .CP(clock), .Q(i[24]) );
  CFD1XL \i_reg[28]  ( .D(n926), .CP(clock), .Q(i[28]) );
  CFD1XL \i_reg[31]  ( .D(n955), .CP(clock), .Q(i[31]) );
  CFD1XL \i_reg[12]  ( .D(n942), .CP(clock), .Q(i[12]), .QN(n2153) );
  CFD1XL \i_reg[2]  ( .D(n950), .CP(clock), .Q(i[2]), .QN(n2156) );
  CFD1XL \i_reg[29]  ( .D(n925), .CP(clock), .Q(i[29]), .QN(n2120) );
  CFD1XL \i_reg[30]  ( .D(n2887), .CP(clock), .Q(i[30]), .QN(n2104) );
  CFD1XL \i_reg[13]  ( .D(n941), .CP(clock), .Q(i[13]), .QN(n2152) );
  CFD1XL \i_reg[14]  ( .D(n940), .CP(clock), .Q(i[14]) );
  CFD1XL \res_not_reg[12]  ( .D(n907), .CP(clock), .Q(res_not_wire[12]), .QN(
        n2147) );
  CFD1XL \result_reg[23]  ( .D(n802), .CP(clock), .Q(result[23]), .QN(n2056)
         );
  CFD1XL \result_reg[26]  ( .D(n2888), .CP(clock), .Q(result[26]), .QN(n2070)
         );
  CFD1XL \result_reg[14]  ( .D(n811), .CP(clock), .Q(result[14]), .QN(n2076)
         );
  CFD1XL \result_reg[27]  ( .D(n2889), .CP(clock), .Q(result[27]), .QN(n2054)
         );
  CFD1XL \result_reg[20]  ( .D(n805), .CP(clock), .Q(result[20]), .QN(n2073)
         );
  CFD1XL \result_reg[17]  ( .D(n808), .CP(clock), .Q(result[17]), .QN(n2059)
         );
  CFD1XL \result_reg[11]  ( .D(n814), .CP(clock), .Q(result[11]), .QN(n2062)
         );
  CFD1XL \result_reg[8]  ( .D(n817), .CP(clock), .Q(result[8]), .QN(n2079) );
  CFD1XL \result_reg[5]  ( .D(n820), .CP(clock), .Q(result[5]), .QN(n2065) );
  CFD1XL \result_reg[2]  ( .D(n823), .CP(clock), .Q(result[2]), .QN(n2081) );
  CFD1XL \result_reg[25]  ( .D(n2890), .CP(clock), .Q(result[25]), .QN(n2055)
         );
  CFD1XL \result_reg[22]  ( .D(n803), .CP(clock), .Q(result[22]), .QN(n2072)
         );
  CFD1XL \result_reg[18]  ( .D(n807), .CP(clock), .Q(result[18]), .QN(n2074)
         );
  CFD1XL \result_reg[16]  ( .D(n809), .CP(clock), .Q(result[16]), .QN(n2075)
         );
  CFD1XL \result_reg[15]  ( .D(n810), .CP(clock), .Q(result[15]), .QN(n2060)
         );
  CFD1XL \result_reg[13]  ( .D(n812), .CP(clock), .Q(result[13]), .QN(n2061)
         );
  CFD1XL \result_reg[12]  ( .D(n2894), .CP(clock), .Q(result[12]), .QN(n2077)
         );
  CFD1XL \result_reg[10]  ( .D(n815), .CP(clock), .Q(result[10]), .QN(n2078)
         );
  CFD1XL \result_reg[9]  ( .D(n2896), .CP(clock), .Q(result[9]), .QN(n2063) );
  CFD1XL \result_reg[7]  ( .D(n818), .CP(clock), .Q(result[7]), .QN(n2064) );
  CFD1XL \result_reg[6]  ( .D(n819), .CP(clock), .Q(result[6]), .QN(n2052) );
  CFD1XL \result_reg[4]  ( .D(n821), .CP(clock), .Q(result[4]), .QN(n2080) );
  CFD1XL \result_reg[3]  ( .D(n822), .CP(clock), .Q(result[3]), .QN(n2066) );
  CFD1XL \result_reg[1]  ( .D(n824), .CP(clock), .Q(result[1]), .QN(n2067) );
  CFD1XL \result_reg[0]  ( .D(n2898), .CP(clock), .Q(result[0]), .QN(n3694) );
  CFD1XL \result_reg[19]  ( .D(n2899), .CP(clock), .Q(result[19]), .QN(n2058)
         );
  CFD1XL \result_reg[24]  ( .D(n2900), .CP(clock), .Q(result[24]), .QN(n2071)
         );
  CFD1XL \result_reg[21]  ( .D(n2901), .CP(clock), .Q(result[21]), .QN(n2057)
         );
  CFD1XL \result_reg[28]  ( .D(n797), .CP(clock), .Q(result[28]), .QN(n2069)
         );
  CFD1XL \res_not_reg[1]  ( .D(n2872), .CP(clock), .QN(n164) );
  CFD1QXL \result_reg[62]  ( .D(n826), .CP(clock), .Q(result[62]) );
  CFD1X1 \result_reg[33]  ( .D(n855), .CP(clock), .Q(result[33]), .QN(n2920)
         );
  CFD1X1 \result_reg[32]  ( .D(n2902), .CP(clock), .Q(result[32]) );
  COND11X1 U1883 ( .A(n3041), .B(i[1]), .C(n2162), .D(n2181), .Z(n951) );
  CENXL U1884 ( .A(n106), .B(n3675), .Z(n3509) );
  CANR1X1 U1885 ( .A(n3535), .B(n3294), .C(n3293), .Z(n3326) );
  CNR2X1 U1886 ( .A(n3605), .B(n3604), .Z(n3394) );
  CENXL U1887 ( .A(n3409), .B(n2091), .Z(n3400) );
  CENXL U1888 ( .A(n3105), .B(n3100), .Z(n3101) );
  CENXL U1889 ( .A(n3095), .B(n3091), .Z(n3092) );
  CENXL U1890 ( .A(n2138), .B(c_inres), .Z(n2634) );
  CENXL U1891 ( .A(n3358), .B(n3357), .Z(n3359) );
  COND2X2 U1892 ( .A(n3332), .B(n2112), .C(n3596), .D(n3595), .Z(n3358) );
  CIVX3 U1893 ( .A(n3116), .Z(n3111) );
  CND2IX2 U1894 ( .B(n3005), .A(n2985), .Z(n3116) );
  CIVX3 U1895 ( .A(n3124), .Z(n3119) );
  CND2X2 U1896 ( .A(n3122), .B(n3057), .Z(n3124) );
  CND2X2 U1897 ( .A(res_not_wire[16]), .B(n3058), .Z(n3102) );
  CENX4 U1898 ( .A(n2957), .B(opera1[31]), .Z(n2956) );
  CND2X2 U1899 ( .A(n3354), .B(n3309), .Z(n3310) );
  CND2X2 U1900 ( .A(n3062), .B(n3061), .Z(n3075) );
  COND3XL U1901 ( .A(n3502), .B(n3501), .C(n3500), .D(n3499), .Z(n826) );
  CANR3X2 U1902 ( .A(n3496), .B(n3661), .C(n3495), .D(n3494), .Z(n3497) );
  CND2X2 U1903 ( .A(n2926), .B(n3063), .Z(n3067) );
  CNR2IX2 U1904 ( .B(res_not_wire[28]), .A(n3071), .Z(n2926) );
  CENXL U1905 ( .A(n3624), .B(n3623), .Z(n3625) );
  COND2X2 U1906 ( .A(n3419), .B(n2036), .C(n3418), .D(n3417), .Z(n3624) );
  CND2X2 U1907 ( .A(n2986), .B(n3454), .Z(n3651) );
  COND1X1 U1908 ( .A(n2956), .B(c_inop1), .C(n3163), .Z(n3514) );
  CND2X1 U1909 ( .A(c_inop1), .B(n2956), .Z(n3163) );
  CND3X2 U1910 ( .A(n2984), .B(res_not_wire[2]), .C(n3157), .Z(n3153) );
  CND2X2 U1911 ( .A(n3053), .B(n3141), .Z(n3143) );
  CAN3XL U1912 ( .A(result[33]), .B(n3165), .C(n3164), .Z(n2862) );
  CND2X2 U1913 ( .A(n3137), .B(n2856), .Z(n3133) );
  CIVX3 U1914 ( .A(n3131), .Z(n3137) );
  CENXL U1915 ( .A(res_not_wire[4]), .B(n3147), .Z(n3148) );
  CND2IX2 U1916 ( .B(n162), .A(n3149), .Z(n3147) );
  CNR3X2 U1917 ( .A(n2103), .B(n2234), .C(n2121), .Z(n2241) );
  CND3X2 U1918 ( .A(i[23]), .B(n2105), .C(i[24]), .Z(n2234) );
  COND1X2 U1919 ( .A(n3046), .B(n2246), .C(i[31]), .Z(n3048) );
  CND3X1 U1920 ( .A(i[27]), .B(n2241), .C(i[28]), .Z(n2246) );
  CIVDX2 U1921 ( .A(n3007), .Z0(n2847), .Z1(n2848) );
  CIVDX2 U1922 ( .A(n3666), .Z0(n2849), .Z1(n2850) );
  CIVDX1 U1923 ( .A(n3008), .Z0(n2851), .Z1(n2852) );
  CND2IXL U1924 ( .B(n3064), .A(n3668), .Z(n3007) );
  CND2IXL U1925 ( .B(n3064), .A(n3010), .Z(n3666) );
  CND2IX1 U1926 ( .B(n3064), .A(n3014), .Z(n3008) );
  CIVXL U1927 ( .A(n2206), .Z(n2145) );
  CND2X2 U1928 ( .A(i[14]), .B(n2206), .Z(n2207) );
  CNR3X2 U1929 ( .A(n2153), .B(n2200), .C(n2152), .Z(n2206) );
  CIVXL U1930 ( .A(n3012), .Z(n2853) );
  CIVXL U1931 ( .A(n3012), .Z(n2854) );
  CDLY1X2 U1932 ( .A(n3668), .Z(n3011) );
  CDLY1X2 U1933 ( .A(n3668), .Z(n3018) );
  CDLY1X2 U1934 ( .A(n3668), .Z(n3017) );
  CDLY1X2 U1935 ( .A(n3668), .Z(n3016) );
  CDLY1X2 U1936 ( .A(n3668), .Z(n3015) );
  CNIVX1 U1937 ( .A(n3668), .Z(n3012) );
  CND2X1 U1938 ( .A(n3462), .B(n3461), .Z(n3476) );
  CND2X1 U1939 ( .A(n3367), .B(n3366), .Z(n3389) );
  CND2X1 U1940 ( .A(n3437), .B(n3436), .Z(n3474) );
  CND2X1 U1941 ( .A(n3493), .B(n3470), .Z(n3491) );
  CND2X1 U1942 ( .A(n3413), .B(n3412), .Z(n3431) );
  CND2X1 U1943 ( .A(n3372), .B(n3371), .Z(n3421) );
  CND2X1 U1944 ( .A(n3272), .B(n3271), .Z(n3282) );
  CND2X1 U1945 ( .A(n3312), .B(n3311), .Z(n3325) );
  CND2X1 U1946 ( .A(n3464), .B(n3463), .Z(n3485) );
  CND2X1 U1947 ( .A(n3316), .B(n3315), .Z(n3337) );
  CND2X1 U1948 ( .A(n3288), .B(n3287), .Z(n3298) );
  CND2X1 U1949 ( .A(n3476), .B(n3475), .Z(n3480) );
  CND2X1 U1950 ( .A(n3389), .B(n3383), .Z(n3384) );
  CND2IX1 U1951 ( .B(n3357), .A(n3358), .Z(n3379) );
  CEOX1 U1952 ( .A(result[61]), .B(n3491), .Z(n3671) );
  CEOX1 U1953 ( .A(result[60]), .B(n3488), .Z(n3503) );
  CEOX1 U1954 ( .A(result[57]), .B(n3479), .Z(n3478) );
  CEOX1 U1955 ( .A(result[58]), .B(n3480), .Z(n3652) );
  CEOX1 U1956 ( .A(result[55]), .B(n3427), .Z(n3633) );
  CEOX1 U1957 ( .A(result[52]), .B(n3395), .Z(n3402) );
  CEOX1 U1958 ( .A(result[47]), .B(n3332), .Z(n3595) );
  CEOX1 U1959 ( .A(result[53]), .B(n3419), .Z(n3418) );
  CND2X1 U1960 ( .A(n3468), .B(n3467), .Z(n3493) );
  CEOX1 U1961 ( .A(result[38]), .B(n3238), .Z(n3576) );
  CEOX1 U1962 ( .A(result[50]), .B(n3384), .Z(n3612) );
  CND2X1 U1963 ( .A(n3411), .B(n3410), .Z(n3423) );
  CND2X1 U1964 ( .A(n3274), .B(n3273), .Z(n3290) );
  CND2X1 U1965 ( .A(n3370), .B(n3369), .Z(n3377) );
  CND2X1 U1966 ( .A(n3314), .B(n3313), .Z(n3321) );
  CND2X1 U1967 ( .A(n3246), .B(n3245), .Z(n3280) );
  CND2X1 U1968 ( .A(n3230), .B(n3229), .Z(n3242) );
  CND3XL U1969 ( .A(n3202), .B(n3201), .C(n3200), .Z(n3236) );
  CND2X1 U1970 ( .A(n3335), .B(n3334), .Z(n3382) );
  CND2X1 U1971 ( .A(n3296), .B(n3295), .Z(n3323) );
  CND2X1 U1972 ( .A(n3429), .B(n3428), .Z(n3439) );
  CND2X1 U1973 ( .A(n3391), .B(n3390), .Z(n3392) );
  CND2X1 U1974 ( .A(n3466), .B(n3465), .Z(n3487) );
  CIVX2 U1975 ( .A(opera2[0]), .Z(n2936) );
  CNIVXL U1976 ( .A(n2643), .Z(n2918) );
  CENX1 U1977 ( .A(opera2[2]), .B(opera2_63), .Z(n2649) );
  CENX1 U1978 ( .A(opera2[25]), .B(opera2_63), .Z(n2795) );
  CANR1X1 U1979 ( .A(n3482), .B(n2928), .C(n3481), .Z(n3641) );
  CEOX1 U1980 ( .A(result[59]), .B(n3483), .Z(n3640) );
  CANR2X1 U1981 ( .A(n3387), .B(n3386), .C(result[50]), .D(n3385), .Z(n3605)
         );
  CANR1XL U1982 ( .A(n3614), .B(n3613), .C(n3612), .Z(n3386) );
  CND3XL U1983 ( .A(n3380), .B(n3614), .C(n3379), .Z(n3387) );
  CEOX1 U1984 ( .A(result[51]), .B(n3392), .Z(n3604) );
  CND2X1 U1985 ( .A(n3194), .B(n3172), .Z(n3191) );
  CEOX1 U1986 ( .A(result[48]), .B(n3333), .Z(n3357) );
  COND1X1 U1987 ( .A(n2862), .B(n3167), .C(n3166), .Z(n3182) );
  CND3X1 U1988 ( .A(i[10]), .B(n2146), .C(i[11]), .Z(n2200) );
  CNR3XL U1989 ( .A(n2157), .B(n2162), .C(n2156), .Z(n2173) );
  CND3XL U1990 ( .A(i[4]), .B(n2150), .C(i[5]), .Z(n2185) );
  CND2X1 U1991 ( .A(i[3]), .B(n2173), .Z(n2180) );
  CND3XL U1992 ( .A(i[8]), .B(n2148), .C(i[9]), .Z(n2195) );
  CND3XL U1993 ( .A(i[15]), .B(n2144), .C(i[16]), .Z(n2212) );
  CND3XL U1994 ( .A(i[17]), .B(n2130), .C(i[18]), .Z(n2217) );
  CND3XL U1995 ( .A(i[19]), .B(n2118), .C(i[20]), .Z(n2222) );
  CND3XL U1996 ( .A(i[21]), .B(n2117), .C(i[22]), .Z(n2227) );
  CENX1 U1997 ( .A(n3448), .B(n3447), .Z(n3449) );
  CENX1 U1998 ( .A(n3653), .B(n3652), .Z(n3654) );
  CEOX1 U1999 ( .A(result[35]), .B(n3191), .Z(n3193) );
  CND3XL U2000 ( .A(i[6]), .B(n2149), .C(i[7]), .Z(n2190) );
  CANR1XL U2001 ( .A(n3261), .B(n3263), .C(n3262), .Z(n3259) );
  CND3XL U2002 ( .A(n3261), .B(n3257), .C(n2948), .Z(n3258) );
  CANR1XL U2003 ( .A(n3567), .B(n3577), .C(n3566), .Z(n3568) );
  CANR1XL U2004 ( .A(n3089), .B(n3088), .C(n3087), .Z(n2778) );
  CNIVX2 U2005 ( .A(n957), .Z(n2884) );
  CENX1 U2006 ( .A(n2989), .B(n3702), .Z(n3445) );
  CND3XL U2007 ( .A(n3639), .B(n3638), .C(n3637), .Z(n834) );
  CENX1 U2008 ( .A(n2983), .B(n3401), .Z(n3408) );
  CND3XL U2009 ( .A(n3560), .B(n3559), .C(n3558), .Z(n846) );
  CENX1 U2010 ( .A(res_not_wire[46]), .B(n3003), .Z(n3601) );
  CENX1 U2011 ( .A(n1053), .B(n3659), .Z(n3667) );
  CENX1 U2012 ( .A(n116), .B(n3611), .Z(n3622) );
  CND2X1 U2013 ( .A(n2802), .B(n2807), .Z(n2813) );
  CAN2X1 U2014 ( .A(res_not_wire[8]), .B(n2863), .Z(n2856) );
  COAN1X1 U2015 ( .A(n2250), .B(n2101), .C(n3047), .Z(n2857) );
  CAN2X1 U2016 ( .A(res_not_wire[20]), .B(n2868), .Z(n2858) );
  CIVDX1 U2017 ( .A(opera1[31]), .Z0(n2859), .Z1(n2860) );
  COR2X1 U2018 ( .A(n2662), .B(n2668), .Z(n2861) );
  CAN2X1 U2019 ( .A(n2722), .B(n3688), .Z(n2864) );
  CEOX1 U2020 ( .A(opera1[5]), .B(opera1[31]), .Z(n2865) );
  COR2X1 U2021 ( .A(n2744), .B(n2738), .Z(n2866) );
  CND2X1 U2022 ( .A(n2944), .B(n2945), .Z(n2635) );
  CNIVX1 U2023 ( .A(n2873), .Z(n2872) );
  CNIVX1 U2024 ( .A(n918), .Z(n2873) );
  CIVXL U2025 ( .A(opera2[30]), .Z(n2003) );
  CIVDX1 U2026 ( .A(n2939), .Z1(n2875) );
  CIVXL U2027 ( .A(opera2[31]), .Z(n2939) );
  CENXL U2028 ( .A(n2875), .B(n2833), .Z(n2829) );
  CND2IXL U2029 ( .B(n3522), .A(n3521), .Z(n794) );
  CNIVX1 U2030 ( .A(n796), .Z(n2876) );
  CEOXL U2031 ( .A(opera2[29]), .B(n2881), .Z(n2820) );
  CNIVX1 U2032 ( .A(n795), .Z(n2877) );
  CDLY1XL U2033 ( .A(start), .Z(n2878) );
  CNR2IXL U2034 ( .B(nst[2]), .A(n2878), .Z(N34) );
  CNIVX1 U2035 ( .A(n2880), .Z(n2879) );
  CNIVX1 U2036 ( .A(n956), .Z(n2880) );
  CNIVXL U2037 ( .A(muordi), .Z(n2885) );
  CNR2XL U2038 ( .A(n2140), .B(n2883), .Z(n2167) );
  CIVX2 U2039 ( .A(opera2_63), .Z(n2002) );
  CNIVX1 U2040 ( .A(n2002), .Z(n2881) );
  CNIVX1 U2041 ( .A(n922), .Z(n2882) );
  CNIVX1 U2042 ( .A(n2885), .Z(n2883) );
  CNIVX1 U2043 ( .A(n928), .Z(n2886) );
  CNIVX1 U2044 ( .A(n924), .Z(n2887) );
  CNIVX1 U2045 ( .A(n799), .Z(n2888) );
  CNIVX1 U2046 ( .A(n798), .Z(n2889) );
  CEOXL U2047 ( .A(opera2[27]), .B(opera2_63), .Z(n2807) );
  CNIVX1 U2048 ( .A(n800), .Z(n2890) );
  CENX1 U2049 ( .A(opera2[22]), .B(opera2_63), .Z(n2776) );
  CNIVX1 U2050 ( .A(n2776), .Z(n2891) );
  CEOXL U2051 ( .A(opera2[18]), .B(opera2_63), .Z(n2750) );
  CENX1 U2052 ( .A(opera2[16]), .B(opera2_63), .Z(n2738) );
  CNIVX1 U2053 ( .A(n2738), .Z(n2892) );
  CEOXL U2054 ( .A(n2737), .B(n2892), .Z(n2734) );
  CEOXL U2055 ( .A(opera2[15]), .B(opera2_63), .Z(n2731) );
  CENX1 U2056 ( .A(opera2[13]), .B(opera2_63), .Z(n2719) );
  CNIVX1 U2057 ( .A(n2719), .Z(n2893) );
  CNIVX1 U2058 ( .A(n813), .Z(n2894) );
  CEOXL U2059 ( .A(opera2[12]), .B(opera2_63), .Z(n2712) );
  CENX1 U2060 ( .A(opera2[10]), .B(opera2_63), .Z(n2700) );
  CNIVX1 U2061 ( .A(n2700), .Z(n2895) );
  CNIVX1 U2062 ( .A(n816), .Z(n2896) );
  CEOXL U2063 ( .A(opera2[9]), .B(opera2_63), .Z(n2693) );
  CENXL U2064 ( .A(opera2[7]), .B(opera2_63), .Z(n2681) );
  CEOXL U2065 ( .A(opera2[6]), .B(opera2_63), .Z(n2674) );
  CENX1 U2066 ( .A(opera2[4]), .B(opera2_63), .Z(n2662) );
  CNIVX1 U2067 ( .A(n2662), .Z(n2897) );
  CEOXL U2068 ( .A(opera2[3]), .B(opera2_63), .Z(n2655) );
  CENXL U2069 ( .A(opera2[1]), .B(opera2_63), .Z(n2642) );
  CNIVX1 U2070 ( .A(n825), .Z(n2898) );
  CNIVX1 U2071 ( .A(n806), .Z(n2899) );
  CENXL U2072 ( .A(opera2[19]), .B(opera2_63), .Z(n2757) );
  CNIVX1 U2073 ( .A(n801), .Z(n2900) );
  CEOXL U2074 ( .A(opera2[24]), .B(opera2_63), .Z(n2788) );
  CNIVX1 U2075 ( .A(n804), .Z(n2901) );
  CEOXL U2076 ( .A(opera2[21]), .B(opera2_63), .Z(n2769) );
  CNIVX1 U2077 ( .A(n856), .Z(n2902) );
  CENX1 U2078 ( .A(opera2[28]), .B(opera2_63), .Z(n2814) );
  CNIVX1 U2079 ( .A(n2814), .Z(n2903) );
  CNR3X1 U2080 ( .A(n2820), .B(n2814), .C(n2813), .Z(n2821) );
  COND1XL U2081 ( .A(n2848), .B(n3512), .C(n3511), .Z(n919) );
  CANR1X1 U2082 ( .A(n3545), .B(n3285), .C(n3284), .Z(n3555) );
  CNR3X2 U2083 ( .A(n2643), .B(n2642), .C(n2649), .Z(n2650) );
  CND2IX1 U2084 ( .B(n3067), .A(n2919), .Z(n3222) );
  CNR2X1 U2085 ( .A(n2993), .B(n2931), .Z(n2919) );
  CANR1XL U2086 ( .A(n3535), .B(n3294), .C(n3293), .Z(n2921) );
  CENX1 U2087 ( .A(opera1[5]), .B(opera1[31]), .Z(n3197) );
  COND2X1 U2088 ( .A(n3286), .B(n2046), .C(n3555), .D(n3554), .Z(n3535) );
  CEOX2 U2089 ( .A(opera1[31]), .B(opera1[1]), .Z(n2922) );
  CNR2X1 U2090 ( .A(n3194), .B(n3199), .Z(n2923) );
  CANR11XL U2091 ( .A(n2847), .B(n3675), .C(n3644), .D(n3643), .Z(n3647) );
  CNR2IX1 U2092 ( .B(res_not_wire[42]), .A(n3551), .Z(n2954) );
  CND3XL U2093 ( .A(res_not_wire[44]), .B(n2954), .C(n3533), .Z(n3344) );
  CIVX2 U2094 ( .A(n3677), .Z(n3659) );
  CNR2X1 U2095 ( .A(n3524), .B(n2953), .Z(n2952) );
  CND2XL U2096 ( .A(n2927), .B(n3190), .Z(n3524) );
  CAN2X1 U2097 ( .A(n3401), .B(n2933), .Z(n2924) );
  CND2IX2 U2098 ( .B(n3611), .A(n2924), .Z(n3409) );
  CNR2IX2 U2099 ( .B(n3091), .A(n3095), .Z(n2925) );
  CNR2IXL U2100 ( .B(n3091), .A(n3095), .Z(n2949) );
  CAN2X2 U2101 ( .A(n2935), .B(n2964), .Z(n3003) );
  CND2X1 U2102 ( .A(n2936), .B(opera2_63), .Z(n2945) );
  CNR2IXL U2103 ( .B(res_not_wire[28]), .A(n3071), .Z(n3001) );
  CNR2IXL U2104 ( .B(n2965), .A(n3222), .Z(n2927) );
  COND2X1 U2105 ( .A(n3479), .B(n2033), .C(n3478), .D(n3477), .Z(n2928) );
  COND2XL U2106 ( .A(n3479), .B(n2033), .C(n3478), .D(n3477), .Z(n3653) );
  COND2XL U2107 ( .A(n3328), .B(n2113), .C(n3327), .D(n2921), .Z(n2929) );
  CNR3X2 U2108 ( .A(n2687), .B(n2681), .C(n2680), .Z(n2688) );
  CNR2X2 U2109 ( .A(n2661), .B(n2861), .Z(n2669) );
  CND2X2 U2110 ( .A(n2991), .B(n2858), .Z(n3095) );
  CND2X1 U2111 ( .A(n2869), .B(res_not_wire[32]), .Z(n2931) );
  CNR2IX2 U2112 ( .B(n2965), .A(n3222), .Z(n2964) );
  CNR3X1 U2113 ( .A(n2706), .B(n2700), .C(n2699), .Z(n2707) );
  CNR2X2 U2114 ( .A(n2737), .B(n2866), .Z(n2745) );
  CNR3X1 U2115 ( .A(n2725), .B(n2719), .C(n2718), .Z(n2726) );
  COND1XL U2116 ( .A(n3588), .B(n3586), .C(n2958), .Z(n3263) );
  CND2IX1 U2117 ( .B(n3389), .A(n3368), .Z(n3391) );
  COR2X1 U2118 ( .A(n3171), .B(n3198), .Z(n3194) );
  CANR4CXL U2119 ( .A(n2738), .B(n2737), .C(n2744), .D(n2745), .Z(n2741) );
  CENX1 U2120 ( .A(n3535), .B(n3534), .Z(n3536) );
  CND2X1 U2121 ( .A(n2669), .B(n2674), .Z(n2680) );
  CENX1 U2122 ( .A(opera1[7]), .B(opera1[31]), .Z(n3239) );
  CENX1 U2123 ( .A(opera1[8]), .B(opera1[31]), .Z(n3233) );
  CENX1 U2124 ( .A(opera1[9]), .B(opera1[31]), .Z(n3247) );
  CEOX1 U2125 ( .A(result[49]), .B(n3378), .Z(n3613) );
  CND3XL U2126 ( .A(n3680), .B(n3679), .C(n3678), .Z(n828) );
  CIVX2 U2127 ( .A(opera2[11]), .Z(n2940) );
  CEOXL U2128 ( .A(opera2[8]), .B(n2002), .Z(n2687) );
  CND3XL U2129 ( .A(n3550), .B(n3549), .C(n3548), .Z(n847) );
  CND3XL U2130 ( .A(n3610), .B(n3609), .C(n3608), .Z(n838) );
  COAN1X1 U2131 ( .A(n2950), .B(n3191), .C(n2951), .Z(n3525) );
  CENX1 U2132 ( .A(opera1[10]), .B(opera1[31]), .Z(n3279) );
  CENX1 U2133 ( .A(opera1[11]), .B(n2860), .Z(n3275) );
  CENX1 U2134 ( .A(opera1[12]), .B(opera1[31]), .Z(n3289) );
  CENX1 U2135 ( .A(opera1[13]), .B(opera1[31]), .Z(n3297) );
  CENX1 U2136 ( .A(opera1[14]), .B(opera1[31]), .Z(n3322) );
  CEOXL U2137 ( .A(opera2[14]), .B(n2002), .Z(n2725) );
  CENX1 U2138 ( .A(opera1[15]), .B(opera1[31]), .Z(n3319) );
  CENX1 U2139 ( .A(opera1[16]), .B(opera1[31]), .Z(n3317) );
  CENX1 U2140 ( .A(opera1[17]), .B(opera1[31]), .Z(n3336) );
  CENX1 U2141 ( .A(opera1[23]), .B(opera1[31]), .Z(n3414) );
  CEOXL U2142 ( .A(opera2[5]), .B(n2002), .Z(n2668) );
  CND2IX2 U2143 ( .B(n2932), .A(c_inres), .Z(n3158) );
  CNR2X1 U2144 ( .A(n3696), .B(n116), .Z(n2933) );
  CIVX2 U2145 ( .A(n3190), .Z(n2934) );
  CNR2X1 U2146 ( .A(n3004), .B(n2934), .Z(n2935) );
  CND2X1 U2147 ( .A(n2650), .B(n2655), .Z(n2661) );
  CANR4CXL U2148 ( .A(n2814), .B(n2813), .C(n2820), .D(n2821), .Z(n2817) );
  CND2XL U2149 ( .A(n2707), .B(n2712), .Z(n2718) );
  CND2XL U2150 ( .A(n2688), .B(n2693), .Z(n2699) );
  CENXL U2151 ( .A(n2826), .B(n2821), .Z(n2824) );
  CND2XL U2152 ( .A(n2764), .B(n2769), .Z(n2775) );
  CND2XL U2153 ( .A(n2783), .B(n2788), .Z(n2794) );
  CEOXL U2154 ( .A(n2813), .B(n2903), .Z(n2810) );
  CEOXL U2155 ( .A(n2794), .B(n2795), .Z(n2791) );
  CEOXL U2156 ( .A(n2775), .B(n2891), .Z(n2772) );
  CND2X1 U2157 ( .A(n3280), .B(n3249), .Z(n3251) );
  CND2X1 U2158 ( .A(n3248), .B(n3234), .Z(n3244) );
  CNR2XL U2159 ( .A(n3488), .B(n2029), .Z(n3489) );
  CNR2XL U2160 ( .A(n3433), .B(n2093), .Z(n3434) );
  CIVX1 U2161 ( .A(n3447), .Z(n3435) );
  CEOXL U2162 ( .A(n2769), .B(n2764), .Z(n2767) );
  CANR1XL U2163 ( .A(n3565), .B(n3576), .C(n3561), .Z(n3588) );
  CND2X1 U2164 ( .A(n3242), .B(n3241), .Z(n3243) );
  CND2X1 U2165 ( .A(n3240), .B(n3239), .Z(n3241) );
  CND2X1 U2166 ( .A(n3282), .B(n3281), .Z(n3283) );
  CND2X1 U2167 ( .A(n3298), .B(n3291), .Z(n3292) );
  CND2X1 U2168 ( .A(n3423), .B(n3422), .Z(n3424) );
  CND2X1 U2169 ( .A(n3325), .B(n3324), .Z(n3329) );
  CEOXL U2170 ( .A(n2731), .B(n2726), .Z(n2729) );
  CND2XL U2171 ( .A(n2952), .B(n3270), .Z(n3541) );
  CEOXL U2172 ( .A(n3612), .B(n2937), .Z(n3618) );
  CANR1XL U2173 ( .A(n3617), .B(n3616), .C(n3615), .Z(n2937) );
  CAN2X1 U2174 ( .A(n3642), .B(n2946), .Z(n3643) );
  CANR4CXL U2175 ( .A(n2719), .B(n2718), .C(n2725), .D(n2726), .Z(n2722) );
  CEOXL U2176 ( .A(n2712), .B(n2707), .Z(n2710) );
  CIVX2 U2177 ( .A(n3673), .Z(n3642) );
  CANR4CXL U2178 ( .A(n2700), .B(n2699), .C(n2706), .D(n2707), .Z(n2703) );
  CNR3XL U2179 ( .A(n2250), .B(n2857), .C(n2137), .Z(n2259) );
  CANR4CXL U2180 ( .A(n2681), .B(n2680), .C(n2687), .D(n2688), .Z(n2684) );
  CEOXL U2181 ( .A(n3561), .B(n3568), .Z(n3569) );
  CND2X1 U2182 ( .A(n2745), .B(n2750), .Z(n2756) );
  CND2XL U2183 ( .A(n2815), .B(n2816), .Z(n796) );
  CND2IX1 U2184 ( .B(n2938), .A(n2823), .Z(n795) );
  CAOR2X2 U2185 ( .A(n3689), .B(result[31]), .C(result[30]), .D(n2854), .Z(
        n2938) );
  CND2XL U2186 ( .A(n2808), .B(n2809), .Z(n797) );
  CND2XL U2187 ( .A(n2796), .B(n2797), .Z(n799) );
  CND2XL U2188 ( .A(n2777), .B(n2778), .Z(n802) );
  CENX1 U2189 ( .A(n2940), .B(n2002), .Z(n2706) );
  CND2IX1 U2190 ( .B(n2941), .A(n2785), .Z(n801) );
  CAOR2X2 U2191 ( .A(n3689), .B(result[25]), .C(result[24]), .D(n2854), .Z(
        n2941) );
  COR2XL U2192 ( .A(n2960), .B(n3238), .Z(n3565) );
  COR2XL U2193 ( .A(n2963), .B(n3243), .Z(n3256) );
  COR2XL U2194 ( .A(n2955), .B(n3244), .Z(n3261) );
  CND2IX1 U2195 ( .B(n2942), .A(n2766), .Z(n804) );
  CAOR2X2 U2196 ( .A(n3689), .B(result[22]), .C(result[21]), .D(n2853), .Z(
        n2942) );
  CND2XL U2197 ( .A(n2751), .B(n2752), .Z(n806) );
  CENX1 U2198 ( .A(n2943), .B(n3493), .Z(n3660) );
  CENX1 U2199 ( .A(result[62]), .B(n3460), .Z(n2943) );
  CIVX8 U2200 ( .A(opera1[0]), .Z(n2957) );
  CND2XL U2201 ( .A(result[34]), .B(n2853), .Z(n2347) );
  COR2XL U2202 ( .A(n2961), .B(n3378), .Z(n3614) );
  CND2IX2 U2203 ( .B(n138), .A(n3073), .Z(n3071) );
  CENXL U2204 ( .A(n2998), .B(n3446), .Z(n3453) );
  COND3X1 U2205 ( .A(n3594), .B(n2852), .C(n3593), .D(n3592), .Z(n849) );
  COND3XL U2206 ( .A(n3543), .B(n3542), .C(n2847), .D(n3551), .Z(n3550) );
  COR2XL U2207 ( .A(n2962), .B(n3333), .Z(n3380) );
  CND2IXL U2208 ( .B(res_not_wire[42]), .A(n3551), .Z(n3552) );
  CIVX1 U2209 ( .A(n160), .Z(n3141) );
  CNR2IXL U2210 ( .B(result[35]), .A(n3011), .Z(n3528) );
  CEOXL U2211 ( .A(n2661), .B(n2897), .Z(n2658) );
  CEOXL U2212 ( .A(n2699), .B(n2895), .Z(n2696) );
  CEOXL U2213 ( .A(n2642), .B(n2918), .Z(n2639) );
  CEOXL U2214 ( .A(n2680), .B(n2681), .Z(n2677) );
  CEOXL U2215 ( .A(n2693), .B(n2688), .Z(n2691) );
  CEOXL U2216 ( .A(n2718), .B(n2893), .Z(n2715) );
  CANR2XL U2217 ( .A(result[34]), .B(n3029), .C(n3023), .D(n2047), .Z(n2297)
         );
  CANR2XL U2218 ( .A(result[35]), .B(n3029), .C(n3023), .D(n2950), .Z(n2298)
         );
  CNR2IXL U2219 ( .B(result[32]), .A(n3013), .Z(n3220) );
  CNR2IXL U2220 ( .B(result[33]), .A(n3017), .Z(n3185) );
  CMXI2XL U2221 ( .A0(n3026), .A1(n3032), .S(result[33]), .Z(n3683) );
  CMXI2XL U2222 ( .A0(n3026), .A1(n3032), .S(result[32]), .Z(n3685) );
  CIVXL U2223 ( .A(result[34]), .Z(n2047) );
  CIVXL U2224 ( .A(res_not_wire[6]), .Z(n2023) );
  CEOXL U2225 ( .A(n2750), .B(n2745), .Z(n2748) );
  CND2X1 U2226 ( .A(opera2[0]), .B(n2002), .Z(n2944) );
  CND2X2 U2227 ( .A(c_inop2), .B(n2635), .Z(n2643) );
  CEOXL U2228 ( .A(c_inop2), .B(n2635), .Z(n2633) );
  CIVX2 U2229 ( .A(n3086), .Z(n3688) );
  CNIVX1 U2230 ( .A(n2179), .Z(n3042) );
  CNIVX1 U2231 ( .A(n2179), .Z(n3043) );
  CIVX2 U2232 ( .A(n2857), .Z(n3034) );
  CNIVX1 U2233 ( .A(n2179), .Z(n3041) );
  CIVX2 U2234 ( .A(n2857), .Z(n3039) );
  CIVX2 U2235 ( .A(n2857), .Z(n3037) );
  CIVX2 U2236 ( .A(n2857), .Z(n3038) );
  CIVX2 U2237 ( .A(n2330), .Z(n3669) );
  CNIVX1 U2238 ( .A(n3668), .Z(n3020) );
  CNIVXL U2239 ( .A(n3668), .Z(n3010) );
  CNIVXL U2240 ( .A(n3668), .Z(n3013) );
  CNIVXL U2241 ( .A(n3668), .Z(n3014) );
  CNIVXL U2242 ( .A(n3668), .Z(n3019) );
  CIVX2 U2243 ( .A(n3075), .Z(n3073) );
  CND2X1 U2244 ( .A(n2857), .B(n2247), .Z(n2178) );
  CND2X1 U2245 ( .A(n3701), .B(n2178), .Z(n2179) );
  CNIVX1 U2246 ( .A(n2259), .Z(n3026) );
  COND1XL U2247 ( .A(n2149), .B(n3043), .C(n2178), .Z(n2187) );
  COND1XL U2248 ( .A(n2146), .B(n3042), .C(n2178), .Z(n2197) );
  COND1XL U2249 ( .A(n2150), .B(n3042), .C(n2178), .Z(n2177) );
  COND1XL U2250 ( .A(n2148), .B(n3043), .C(n2178), .Z(n2192) );
  COND1XL U2251 ( .A(n2144), .B(n3042), .C(n2178), .Z(n2209) );
  COND1XL U2252 ( .A(n2118), .B(n3042), .C(n2178), .Z(n2219) );
  COND1XL U2253 ( .A(n2130), .B(n3042), .C(n2178), .Z(n2214) );
  COND1XL U2254 ( .A(n2117), .B(n3042), .C(n2178), .Z(n2224) );
  COND1XL U2255 ( .A(n2105), .B(n3042), .C(n2178), .Z(n2229) );
  CNIVX1 U2256 ( .A(n2259), .Z(n3023) );
  CNIVX1 U2257 ( .A(n2259), .Z(n3024) );
  CNIVX1 U2258 ( .A(n2259), .Z(n3025) );
  CNIVX1 U2259 ( .A(n2259), .Z(n3022) );
  CNIVX1 U2260 ( .A(n2259), .Z(n3021) );
  CAN2X1 U2261 ( .A(n2247), .B(n2140), .Z(n2249) );
  CNR3XL U2262 ( .A(n2763), .B(n2757), .C(n2756), .Z(n2764) );
  CNR3XL U2263 ( .A(n2801), .B(n2795), .C(n2794), .Z(n2802) );
  CNR3XL U2264 ( .A(n2782), .B(n2776), .C(n2775), .Z(n2783) );
  CND2X1 U2265 ( .A(n3694), .B(n3689), .Z(n2330) );
  CANR1XL U2266 ( .A(n3194), .B(n3199), .C(n2923), .Z(n3195) );
  CENX1 U2267 ( .A(n3000), .B(n2116), .Z(n3175) );
  CNR2XL U2268 ( .A(n3480), .B(n2034), .Z(n3481) );
  CND2X1 U2269 ( .A(n2726), .B(n2731), .Z(n2737) );
  CNR2X1 U2270 ( .A(n3329), .B(n2040), .Z(n3330) );
  CNR2X1 U2271 ( .A(n3283), .B(n2044), .Z(n3284) );
  CND2IX1 U2272 ( .B(n3564), .A(n3526), .Z(n3254) );
  CEOXL U2273 ( .A(n3477), .B(n3478), .Z(n3441) );
  CNR2X1 U2274 ( .A(n3424), .B(n2035), .Z(n3425) );
  CNR2X1 U2275 ( .A(n3292), .B(n2115), .Z(n3293) );
  COND1XL U2276 ( .A(n2923), .B(n2865), .C(n3236), .Z(n3204) );
  CNR2XL U2277 ( .A(n3392), .B(n2097), .Z(n3393) );
  CNR2X1 U2278 ( .A(n3197), .B(n3196), .Z(n3201) );
  CNIVX1 U2279 ( .A(n2927), .Z(n3000) );
  CND2X1 U2280 ( .A(n3277), .B(n3278), .Z(n3545) );
  CENX1 U2281 ( .A(n2881), .B(n2003), .Z(n2826) );
  CND2XL U2282 ( .A(n3487), .B(n3469), .Z(n3470) );
  CND2X1 U2283 ( .A(n3485), .B(n3472), .Z(n3483) );
  CND2XL U2284 ( .A(n3476), .B(n3471), .Z(n3472) );
  CND2X1 U2285 ( .A(n3377), .B(n3376), .Z(n3395) );
  CND2X1 U2286 ( .A(n3391), .B(n3375), .Z(n3376) );
  CND2X1 U2287 ( .A(n3431), .B(n3415), .Z(n3427) );
  CND2XL U2288 ( .A(n3423), .B(n3414), .Z(n3415) );
  CND2X1 U2289 ( .A(n3474), .B(n3440), .Z(n3479) );
  CND2XL U2290 ( .A(n3439), .B(n3438), .Z(n3440) );
  CND2X1 U2291 ( .A(n3421), .B(n3374), .Z(n3419) );
  CND2XL U2292 ( .A(n3377), .B(n3373), .Z(n3374) );
  CND2XL U2293 ( .A(n3321), .B(n3320), .Z(n3332) );
  CND2XL U2294 ( .A(n3325), .B(n3319), .Z(n3320) );
  CND2XL U2295 ( .A(n3290), .B(n3276), .Z(n3286) );
  CND2XL U2296 ( .A(n3282), .B(n3275), .Z(n3276) );
  CNR2IX1 U2297 ( .B(n2779), .A(n3086), .Z(n3087) );
  CND2XL U2298 ( .A(n3280), .B(n3279), .Z(n3281) );
  CND2XL U2299 ( .A(n3290), .B(n3289), .Z(n3291) );
  CND2X1 U2300 ( .A(n3487), .B(n3486), .Z(n3488) );
  CND2XL U2301 ( .A(n3485), .B(n3484), .Z(n3486) );
  CND2XL U2302 ( .A(n3474), .B(n3473), .Z(n3475) );
  CND2XL U2303 ( .A(n3389), .B(n3388), .Z(n3390) );
  CND2XL U2304 ( .A(n3439), .B(n3432), .Z(n3433) );
  CND2XL U2305 ( .A(n3431), .B(n3430), .Z(n3432) );
  CND2XL U2306 ( .A(n3421), .B(n3420), .Z(n3422) );
  CND2XL U2307 ( .A(n3323), .B(n3322), .Z(n3324) );
  CND2XL U2308 ( .A(n3202), .B(n3160), .Z(n3171) );
  CNR2IXL U2309 ( .B(n2849), .A(n2952), .Z(n3208) );
  CNR2IXL U2310 ( .B(n2847), .A(n2954), .Z(n3553) );
  CND2XL U2311 ( .A(n3382), .B(n3381), .Z(n3383) );
  CND2XL U2312 ( .A(n3382), .B(n3338), .Z(n3378) );
  CND2XL U2313 ( .A(n3337), .B(n3336), .Z(n3338) );
  CND2XL U2314 ( .A(n3171), .B(n3198), .Z(n3172) );
  CND2XL U2315 ( .A(n3240), .B(n3237), .Z(n3238) );
  CND2XL U2316 ( .A(n3236), .B(n3235), .Z(n3237) );
  CND2XL U2317 ( .A(n3337), .B(n3318), .Z(n3333) );
  CND2XL U2318 ( .A(n3321), .B(n3317), .Z(n3318) );
  CND2XL U2319 ( .A(n3242), .B(n3233), .Z(n3234) );
  CND2XL U2320 ( .A(n3323), .B(n3299), .Z(n3328) );
  CND2XL U2321 ( .A(n3298), .B(n3297), .Z(n3299) );
  CND3XL U2322 ( .A(n3225), .B(n3224), .C(n3223), .Z(n856) );
  CND2X1 U2323 ( .A(n2252), .B(n3047), .Z(n3050) );
  CND2XL U2324 ( .A(n3162), .B(n3163), .Z(n3164) );
  CEOXL U2325 ( .A(n3641), .B(n3640), .Z(n2946) );
  CNR2IXL U2326 ( .B(n3214), .A(n3673), .Z(n3217) );
  CNIVXL U2327 ( .A(n3630), .Z(n2996) );
  CND3XL U2328 ( .A(n3189), .B(n3188), .C(n3187), .Z(n855) );
  CND2XL U2329 ( .A(n3642), .B(n3184), .Z(n3188) );
  CANR1XL U2330 ( .A(n3186), .B(n3669), .C(n3185), .Z(n3187) );
  CNR2X1 U2331 ( .A(n2051), .B(n3018), .Z(n3519) );
  CNR2IX1 U2332 ( .B(n3078), .A(n3697), .Z(n3062) );
  CNR2IX1 U2333 ( .B(n3523), .A(n2116), .Z(n3190) );
  CND2XL U2334 ( .A(n3248), .B(n3247), .Z(n3249) );
  CND2XL U2335 ( .A(n3165), .B(n3164), .Z(n3215) );
  CND2XL U2336 ( .A(n3171), .B(n3161), .Z(n3168) );
  CND2XL U2337 ( .A(n3165), .B(n3196), .Z(n3161) );
  CNR2XL U2338 ( .A(n2947), .B(n3673), .Z(n3339) );
  CEOX1 U2339 ( .A(n3616), .B(n3613), .Z(n2947) );
  CND2XL U2340 ( .A(n3562), .B(n3565), .Z(n3585) );
  CNR2IX1 U2341 ( .B(n3256), .A(n3585), .Z(n2948) );
  CEOXL U2342 ( .A(n3633), .B(n3634), .Z(n3635) );
  CEOXL U2343 ( .A(n3402), .B(n3403), .Z(n3404) );
  CNIVX1 U2344 ( .A(n2258), .Z(n3029) );
  CNIVX1 U2345 ( .A(n2258), .Z(n3031) );
  CND2XL U2346 ( .A(n3379), .B(n3380), .Z(n3616) );
  CNIVX1 U2347 ( .A(n2258), .Z(n3032) );
  CENX1 U2348 ( .A(n2929), .B(n3345), .Z(n3347) );
  CEOXL U2349 ( .A(n3604), .B(n3605), .Z(n3606) );
  CANR1XL U2350 ( .A(n2246), .B(n3044), .C(n2007), .Z(n2242) );
  CANR1XL U2351 ( .A(n2234), .B(n3044), .C(n2007), .Z(n2232) );
  CANR1XL U2352 ( .A(n2157), .B(n3044), .C(n2182), .Z(n2170) );
  CANR1XL U2353 ( .A(n2834), .B(n3691), .C(n2256), .Z(n3047) );
  CNIVX1 U2354 ( .A(n2258), .Z(n3028) );
  CNIVX1 U2355 ( .A(n2258), .Z(n3027) );
  CANR1XL U2356 ( .A(n2200), .B(n3044), .C(n2007), .Z(n2202) );
  CEOXL U2357 ( .A(n3595), .B(n3596), .Z(n3597) );
  COND2X1 U2358 ( .A(n2242), .B(n2120), .C(n3041), .D(n2243), .Z(n925) );
  CND2X1 U2359 ( .A(n3700), .B(n2120), .Z(n2243) );
  COND2X1 U2360 ( .A(n2232), .B(n2103), .C(n3041), .D(n2233), .Z(n929) );
  CEOX1 U2361 ( .A(n2756), .B(n2757), .Z(n2753) );
  CNIVX1 U2362 ( .A(n2258), .Z(n3030) );
  CND2X1 U2363 ( .A(n2837), .B(n3701), .Z(n2247) );
  COND4CX1 U2364 ( .A(n2170), .B(n2171), .C(n2151), .D(n2172), .Z(n954) );
  CANR11XL U2365 ( .A(n2173), .B(n2151), .C(n3044), .D(n2008), .Z(n2172) );
  CND2XL U2366 ( .A(n3044), .B(n2156), .Z(n2171) );
  CEOXL U2367 ( .A(n2921), .B(n3327), .Z(n3300) );
  CEOXL U2368 ( .A(n3554), .B(n3555), .Z(n3556) );
  CENX1 U2369 ( .A(n2958), .B(n3589), .Z(n3590) );
  CANR1XL U2370 ( .A(n3588), .B(n3587), .C(n3586), .Z(n3589) );
  COND3XL U2371 ( .A(n3264), .B(n3263), .C(n3262), .D(n3261), .Z(n3265) );
  CND2X1 U2372 ( .A(n3699), .B(n2141), .Z(n2254) );
  CANR1XL U2373 ( .A(n2255), .B(n3701), .C(n2256), .Z(n2253) );
  CND2XL U2374 ( .A(n3562), .B(n3584), .Z(n3577) );
  CNIVXL U2375 ( .A(n3117), .Z(n2988) );
  CEOXL U2376 ( .A(n3133), .B(n2159), .Z(n3129) );
  CENX1 U2377 ( .A(n2987), .B(n3157), .Z(n3159) );
  CEOXL U2378 ( .A(n3143), .B(n2023), .Z(n3139) );
  CNR3XL U2379 ( .A(n3214), .B(n2250), .C(n3694), .Z(n3218) );
  CNIVXL U2380 ( .A(n3158), .Z(n2987) );
  COR2X1 U2381 ( .A(n3193), .B(n3192), .Z(n2951) );
  CENX1 U2382 ( .A(opera1[6]), .B(opera1[31]), .Z(n3235) );
  CND4X1 U2383 ( .A(res_not_wire[40]), .B(n3270), .C(n2952), .D(n3542), .Z(
        n3551) );
  CEOX1 U2384 ( .A(result[39]), .B(n3243), .Z(n3561) );
  CEOX1 U2385 ( .A(result[43]), .B(n3286), .Z(n3554) );
  CEOX1 U2386 ( .A(result[42]), .B(n3283), .Z(n3544) );
  CNR2IXL U2387 ( .B(result[62]), .A(n3493), .Z(n3495) );
  CANR1XL U2388 ( .A(n3695), .B(n3493), .C(n3492), .Z(n3494) );
  CEOX1 U2389 ( .A(result[45]), .B(n3328), .Z(n3327) );
  CNR2IXL U2390 ( .B(n3513), .A(n3673), .Z(n3517) );
  CND2XL U2391 ( .A(n2330), .B(n3515), .Z(n3516) );
  CND2XL U2392 ( .A(n3689), .B(n3514), .Z(n3515) );
  CEOX1 U2393 ( .A(result[44]), .B(n3292), .Z(n3534) );
  CEOX1 U2394 ( .A(result[56]), .B(n3433), .Z(n3447) );
  CEOX1 U2395 ( .A(result[54]), .B(n3424), .Z(n3623) );
  CEOX1 U2396 ( .A(result[46]), .B(n3329), .Z(n3345) );
  CNR2IX1 U2397 ( .B(res_not_wire[40]), .A(n3541), .Z(n3543) );
  CND2X1 U2398 ( .A(i[30]), .B(i[29]), .Z(n3046) );
  CND3XL U2399 ( .A(n3642), .B(n3278), .C(n3265), .Z(n3268) );
  CANR1XL U2400 ( .A(result[41]), .B(n3669), .C(n3266), .Z(n3267) );
  CANR1XL U2401 ( .A(n3533), .B(n2954), .C(res_not_wire[44]), .Z(n3305) );
  CND2XL U2402 ( .A(n3642), .B(n3300), .Z(n3303) );
  CND2XL U2403 ( .A(n3642), .B(n3396), .Z(n3399) );
  CANR1XL U2404 ( .A(result[53]), .B(n3669), .C(n3397), .Z(n3398) );
  CND2XL U2405 ( .A(n3642), .B(n3441), .Z(n3444) );
  CANR1XL U2406 ( .A(result[57]), .B(n3669), .C(n3442), .Z(n3443) );
  CANR1XL U2407 ( .A(result[60]), .B(n3669), .C(n3506), .Z(n3507) );
  CND2XL U2408 ( .A(n3642), .B(n3527), .Z(n3530) );
  CANR1XL U2409 ( .A(n3575), .B(n2952), .C(res_not_wire[38]), .Z(n3574) );
  CND2XL U2410 ( .A(n3642), .B(n3569), .Z(n3572) );
  CND2XL U2411 ( .A(n3642), .B(n3597), .Z(n3600) );
  CANR1XL U2412 ( .A(result[47]), .B(n3669), .C(n3598), .Z(n3599) );
  CANR1XL U2413 ( .A(result[45]), .B(n3669), .C(n3301), .Z(n3302) );
  CNR2IX1 U2414 ( .B(result[44]), .A(n3015), .Z(n3301) );
  CANR1XL U2415 ( .A(result[36]), .B(n3669), .C(n3528), .Z(n3529) );
  CANR1XL U2416 ( .A(result[39]), .B(n3669), .C(n3570), .Z(n3571) );
  CNR2IX1 U2417 ( .B(result[38]), .A(n3015), .Z(n3570) );
  CND2IX1 U2418 ( .B(n3673), .A(n3498), .Z(n3499) );
  CANR1XL U2419 ( .A(result[62]), .B(n3669), .C(n3663), .Z(n3664) );
  CENX1 U2420 ( .A(result[40]), .B(n3244), .Z(n2958) );
  COND3X1 U2421 ( .A(n3453), .B(n2850), .C(n3452), .D(n3451), .Z(n833) );
  CND2XL U2422 ( .A(n3642), .B(n3449), .Z(n3452) );
  CANR1XL U2423 ( .A(result[56]), .B(n3669), .C(n3450), .Z(n3451) );
  COND3XL U2424 ( .A(n2950), .B(n2330), .C(n2347), .D(n2348), .Z(n854) );
  COND3X1 U2425 ( .A(n3351), .B(n2852), .C(n3350), .D(n3349), .Z(n843) );
  CND2XL U2426 ( .A(n3642), .B(n3347), .Z(n3350) );
  CANR1XL U2427 ( .A(result[46]), .B(n3669), .C(n3348), .Z(n3349) );
  COND3X1 U2428 ( .A(n3408), .B(n2852), .C(n3407), .D(n3406), .Z(n837) );
  CND2XL U2429 ( .A(n3642), .B(n3404), .Z(n3407) );
  CANR1XL U2430 ( .A(result[52]), .B(n3669), .C(n3405), .Z(n3406) );
  COND3X1 U2431 ( .A(n3540), .B(n2848), .C(n3539), .D(n3538), .Z(n845) );
  CND2XL U2432 ( .A(n3642), .B(n3536), .Z(n3539) );
  CANR1XL U2433 ( .A(result[44]), .B(n3669), .C(n3537), .Z(n3538) );
  COND3X1 U2434 ( .A(n3582), .B(n2848), .C(n3581), .D(n3580), .Z(n851) );
  CND2XL U2435 ( .A(n3642), .B(n3578), .Z(n3581) );
  CANR1XL U2436 ( .A(result[38]), .B(n3669), .C(n3579), .Z(n3580) );
  CND2XL U2437 ( .A(n3642), .B(n3590), .Z(n3593) );
  CANR1XL U2438 ( .A(result[40]), .B(n3669), .C(n3591), .Z(n3592) );
  COND3X1 U2439 ( .A(n3622), .B(n2852), .C(n3621), .D(n3620), .Z(n839) );
  CND2XL U2440 ( .A(n3642), .B(n3618), .Z(n3621) );
  CANR1XL U2441 ( .A(result[50]), .B(n3669), .C(n3619), .Z(n3620) );
  CNR2XL U2442 ( .A(n3630), .B(n2959), .Z(n2998) );
  CANR2X1 U2443 ( .A(n2821), .B(n2003), .C(n2001), .D(n2881), .Z(n2833) );
  CNR2IX1 U2444 ( .B(result[61]), .A(n3015), .Z(n3663) );
  CNR2IX1 U2445 ( .B(result[36]), .A(n3011), .Z(n3209) );
  CNR2IX1 U2446 ( .B(result[40]), .A(n3017), .Z(n3266) );
  CNR2IX1 U2447 ( .B(result[48]), .A(n3012), .Z(n3341) );
  CNR2IX1 U2448 ( .B(result[45]), .A(n3017), .Z(n3348) );
  CNR2IX1 U2449 ( .B(result[47]), .A(n3012), .Z(n3360) );
  CNR2IX1 U2450 ( .B(result[52]), .A(n3016), .Z(n3397) );
  CNR2IX1 U2451 ( .B(result[51]), .A(n3011), .Z(n3405) );
  CNR2IX1 U2452 ( .B(result[56]), .A(n3018), .Z(n3442) );
  CNR2IX1 U2453 ( .B(result[55]), .A(n3012), .Z(n3450) );
  CNR2IX1 U2454 ( .B(result[59]), .A(n3015), .Z(n3506) );
  CNR2IX1 U2455 ( .B(result[43]), .A(n3018), .Z(n3537) );
  CNR2IX1 U2456 ( .B(result[41]), .A(n3011), .Z(n3547) );
  CNR2IX1 U2457 ( .B(result[42]), .A(n3016), .Z(n3557) );
  CNR2IX1 U2458 ( .B(result[37]), .A(n3011), .Z(n3579) );
  CNR2IX1 U2459 ( .B(result[39]), .A(n3018), .Z(n3591) );
  CNR2IX1 U2460 ( .B(result[46]), .A(n3017), .Z(n3598) );
  CNR2IX1 U2461 ( .B(result[50]), .A(n3018), .Z(n3607) );
  CNR2IX1 U2462 ( .B(result[49]), .A(n3016), .Z(n3619) );
  CNR2IX1 U2463 ( .B(result[53]), .A(n3017), .Z(n3626) );
  CNR2IX1 U2464 ( .B(result[54]), .A(n3013), .Z(n3636) );
  CNR2IX1 U2465 ( .B(result[57]), .A(n3015), .Z(n3655) );
  CND3XL U2466 ( .A(res_not_wire[38]), .B(n2952), .C(n3575), .Z(n3583) );
  CND2X1 U2467 ( .A(n3277), .B(n3252), .Z(n3262) );
  CND2X1 U2468 ( .A(res_not_wire[42]), .B(res_not_wire[40]), .Z(n3307) );
  CND3XL U2469 ( .A(n3629), .B(n3628), .C(n3627), .Z(n835) );
  CND2XL U2470 ( .A(n3642), .B(n3625), .Z(n3628) );
  CANR1XL U2471 ( .A(result[54]), .B(n3669), .C(n3626), .Z(n3627) );
  CND3XL U2472 ( .A(n3658), .B(n3657), .C(n3656), .Z(n831) );
  CANR1XL U2473 ( .A(result[58]), .B(n3669), .C(n3655), .Z(n3656) );
  CND2X1 U2474 ( .A(result[41]), .B(n3250), .Z(n3277) );
  CANR2XL U2475 ( .A(result[60]), .B(n2853), .C(result[61]), .D(n3669), .Z(
        n3680) );
  CND2XL U2476 ( .A(n3642), .B(n3635), .Z(n3638) );
  CANR1XL U2477 ( .A(result[55]), .B(n3669), .C(n3636), .Z(n3637) );
  CND3XL U2478 ( .A(n3363), .B(n3362), .C(n3361), .Z(n841) );
  CND2XL U2479 ( .A(n3642), .B(n3359), .Z(n3362) );
  CND2X1 U2480 ( .A(n3356), .B(n3355), .Z(n3363) );
  CANR1XL U2481 ( .A(result[48]), .B(n3669), .C(n3360), .Z(n3361) );
  CND2XL U2482 ( .A(n3642), .B(n3546), .Z(n3549) );
  CANR1XL U2483 ( .A(result[42]), .B(n3669), .C(n3547), .Z(n3548) );
  CND2X1 U2484 ( .A(n3553), .B(n3552), .Z(n3560) );
  CND2XL U2485 ( .A(n3642), .B(n3556), .Z(n3559) );
  CANR1XL U2486 ( .A(result[43]), .B(n3669), .C(n3557), .Z(n3558) );
  CND2XL U2487 ( .A(n3642), .B(n3606), .Z(n3609) );
  CND2X1 U2488 ( .A(n3603), .B(n3602), .Z(n3610) );
  CANR1XL U2489 ( .A(result[51]), .B(n3669), .C(n3607), .Z(n3608) );
  CNR2X1 U2490 ( .A(n106), .B(n3674), .Z(n3457) );
  CANR1XL U2491 ( .A(result[59]), .B(n3669), .C(n3645), .Z(n3646) );
  CNR2IX1 U2492 ( .B(result[58]), .A(n3016), .Z(n3645) );
  CANR2XL U2493 ( .A(n3689), .B(result[15]), .C(result[14]), .D(n2853), .Z(
        n2720) );
  CNR2IX1 U2494 ( .B(result[62]), .A(n3016), .Z(n3459) );
  CENX1 U2495 ( .A(n134), .B(n2992), .Z(n3520) );
  CND2X1 U2496 ( .A(n3211), .B(n3210), .Z(n852) );
  CANR2XL U2497 ( .A(n3208), .B(n3207), .C(n3642), .D(n3206), .Z(n3211) );
  CANR1XL U2498 ( .A(result[37]), .B(n3669), .C(n3209), .Z(n3210) );
  CND2X1 U2499 ( .A(n3343), .B(n3342), .Z(n840) );
  CANR1XL U2500 ( .A(result[49]), .B(n3669), .C(n3341), .Z(n3342) );
  CND2X1 U2501 ( .A(n2630), .B(n2631), .Z(n825) );
  CANR2X1 U2502 ( .A(n3688), .B(n2633), .C(n2847), .D(n2634), .Z(n2631) );
  CANR2XL U2503 ( .A(n3689), .B(result[1]), .C(n2853), .D(result[0]), .Z(n2630) );
  CND2X1 U2504 ( .A(n2656), .B(n2657), .Z(n821) );
  CANR2X1 U2505 ( .A(n2658), .B(n3688), .C(n2847), .D(n3148), .Z(n2657) );
  CANR2XL U2506 ( .A(n3689), .B(result[5]), .C(result[4]), .D(n3009), .Z(n2656) );
  CND2X1 U2507 ( .A(n2682), .B(n2683), .Z(n817) );
  CANR2XL U2508 ( .A(n3689), .B(result[9]), .C(result[8]), .D(n2854), .Z(n2682) );
  CND2X1 U2509 ( .A(n2694), .B(n2695), .Z(n815) );
  CANR2X1 U2510 ( .A(n2696), .B(n3688), .C(n2851), .D(n3128), .Z(n2695) );
  CANR2XL U2511 ( .A(n3689), .B(result[11]), .C(result[10]), .D(n2853), .Z(
        n2694) );
  CND2X1 U2512 ( .A(n2708), .B(n2709), .Z(n813) );
  CANR2X1 U2513 ( .A(n2710), .B(n3688), .C(n2851), .D(n3120), .Z(n2709) );
  CANR2XL U2514 ( .A(n3689), .B(result[13]), .C(result[12]), .D(n3009), .Z(
        n2708) );
  CENX1 U2515 ( .A(n2147), .B(n3119), .Z(n3120) );
  CND2X1 U2516 ( .A(n2732), .B(n2733), .Z(n809) );
  CANR2X1 U2517 ( .A(n2734), .B(n3688), .C(n2849), .D(n3110), .Z(n2733) );
  CANR2XL U2518 ( .A(n3689), .B(result[17]), .C(result[16]), .D(n3009), .Z(
        n2732) );
  CENX1 U2519 ( .A(res_not_wire[16]), .B(n3109), .Z(n3110) );
  CND2X1 U2520 ( .A(n2746), .B(n2747), .Z(n807) );
  CANR2X1 U2521 ( .A(n2748), .B(n3688), .C(n2851), .D(n3101), .Z(n2747) );
  CANR2XL U2522 ( .A(n3689), .B(result[19]), .C(result[18]), .D(n3009), .Z(
        n2746) );
  CND2X1 U2523 ( .A(n2758), .B(n2759), .Z(n805) );
  CANR2XL U2524 ( .A(n3689), .B(result[21]), .C(result[20]), .D(n2854), .Z(
        n2758) );
  CND2X1 U2525 ( .A(n2770), .B(n2771), .Z(n803) );
  CANR2X1 U2526 ( .A(n2772), .B(n3688), .C(n2851), .D(n3090), .Z(n2771) );
  CANR2XL U2527 ( .A(n3689), .B(result[23]), .C(result[22]), .D(n2854), .Z(
        n2770) );
  CENX1 U2528 ( .A(n2949), .B(n2126), .Z(n3090) );
  CANR2X1 U2529 ( .A(n2786), .B(n3688), .C(n2847), .D(n3082), .Z(n2785) );
  CENX1 U2530 ( .A(n2124), .B(n3081), .Z(n3082) );
  CANR2XL U2531 ( .A(n3689), .B(result[27]), .C(result[26]), .D(n3009), .Z(
        n2796) );
  CANR2XL U2532 ( .A(n3689), .B(result[29]), .C(result[28]), .D(n3009), .Z(
        n2808) );
  CENX1 U2533 ( .A(res_not_wire[28]), .B(n3071), .Z(n3072) );
  CND2X1 U2534 ( .A(n2637), .B(n2638), .Z(n824) );
  CANR2X1 U2535 ( .A(n2639), .B(n3688), .C(n2851), .D(n3159), .Z(n2638) );
  CANR2XL U2536 ( .A(n3689), .B(result[2]), .C(result[1]), .D(n3009), .Z(n2637) );
  CND2X1 U2537 ( .A(n2651), .B(n2652), .Z(n822) );
  CANR2X1 U2538 ( .A(n2653), .B(n3688), .C(n2851), .D(n3150), .Z(n2652) );
  CANR2XL U2539 ( .A(n3689), .B(result[4]), .C(result[3]), .D(n3009), .Z(n2651) );
  CND2X1 U2540 ( .A(n2663), .B(n2664), .Z(n820) );
  CANR2XL U2541 ( .A(n3689), .B(result[6]), .C(result[5]), .D(n2854), .Z(n2663) );
  CND2X1 U2542 ( .A(n2675), .B(n2676), .Z(n818) );
  CANR2X1 U2543 ( .A(n2677), .B(n3688), .C(n2849), .D(n3138), .Z(n2676) );
  CANR2XL U2544 ( .A(n3689), .B(result[8]), .C(result[7]), .D(n2853), .Z(n2675) );
  CND2X1 U2545 ( .A(n2689), .B(n2690), .Z(n816) );
  CANR2X1 U2546 ( .A(n2691), .B(n3688), .C(n2849), .D(n3129), .Z(n2690) );
  CANR2XL U2547 ( .A(n3689), .B(result[10]), .C(result[9]), .D(n3009), .Z(
        n2689) );
  CND2X1 U2548 ( .A(n2701), .B(n2702), .Z(n814) );
  CANR2XL U2549 ( .A(n3689), .B(result[12]), .C(result[11]), .D(n2854), .Z(
        n2701) );
  CND2X1 U2550 ( .A(n2713), .B(n2714), .Z(n812) );
  CANR2X1 U2551 ( .A(n2715), .B(n3688), .C(n2847), .D(n3118), .Z(n2714) );
  CANR2XL U2552 ( .A(n3689), .B(result[14]), .C(result[13]), .D(n2853), .Z(
        n2713) );
  CND2X1 U2553 ( .A(n2727), .B(n2728), .Z(n810) );
  CANR2X1 U2554 ( .A(n2729), .B(n3688), .C(n2847), .D(n3112), .Z(n2728) );
  CANR2XL U2555 ( .A(n3689), .B(result[16]), .C(result[15]), .D(n3009), .Z(
        n2727) );
  CENX1 U2556 ( .A(n150), .B(n3111), .Z(n3112) );
  CND2X1 U2557 ( .A(n2739), .B(n2740), .Z(n808) );
  CANR2XL U2558 ( .A(n3689), .B(result[18]), .C(result[17]), .D(n2854), .Z(
        n2739) );
  CANR2X1 U2559 ( .A(n2753), .B(n3688), .C(n2847), .D(n3099), .Z(n2752) );
  CANR2XL U2560 ( .A(n3689), .B(result[20]), .C(result[19]), .D(n3009), .Z(
        n2751) );
  CENX1 U2561 ( .A(n146), .B(n2990), .Z(n3099) );
  CANR2XL U2562 ( .A(n3689), .B(result[24]), .C(result[23]), .D(n2854), .Z(
        n2777) );
  CND2X1 U2563 ( .A(n2789), .B(n2790), .Z(n800) );
  CANR2X1 U2564 ( .A(n2791), .B(n3688), .C(n2851), .D(n3080), .Z(n2790) );
  CANR2XL U2565 ( .A(n3689), .B(result[26]), .C(result[25]), .D(n3009), .Z(
        n2789) );
  CENX1 U2566 ( .A(n3079), .B(n3078), .Z(n3080) );
  CND2X1 U2567 ( .A(n2803), .B(n2804), .Z(n798) );
  CANR2XL U2568 ( .A(n3689), .B(result[28]), .C(result[27]), .D(n3009), .Z(
        n2803) );
  CENX1 U2569 ( .A(n138), .B(n3073), .Z(n3074) );
  CANR2XL U2570 ( .A(n3689), .B(result[30]), .C(result[29]), .D(n3009), .Z(
        n2815) );
  CND2X1 U2571 ( .A(n2670), .B(n2671), .Z(n819) );
  CANR2X1 U2572 ( .A(n2672), .B(n3688), .C(n2849), .D(n3139), .Z(n2671) );
  CANR2XL U2573 ( .A(n3689), .B(result[7]), .C(result[6]), .D(n3009), .Z(n2670) );
  CND2X1 U2574 ( .A(n2644), .B(n2645), .Z(n823) );
  CANR2XL U2575 ( .A(n3689), .B(result[3]), .C(result[2]), .D(n2853), .Z(n2644) );
  CND2X1 U2576 ( .A(n2151), .B(n2155), .Z(n2839) );
  COND1XL U2577 ( .A(n3033), .B(n2050), .C(n2838), .Z(n793) );
  COND1XL U2578 ( .A(n3035), .B(n2993), .C(n2293), .Z(n889) );
  CANR2X1 U2579 ( .A(result[30]), .B(n3029), .C(n3023), .D(n2068), .Z(n2293)
         );
  COND1XL U2580 ( .A(n3033), .B(n2090), .C(n2317), .Z(n865) );
  CANR2X1 U2581 ( .A(result[54]), .B(n3031), .C(n3025), .D(n2035), .Z(n2317)
         );
  CND2IX1 U2582 ( .B(i[31]), .A(n2843), .Z(n2837) );
  CNR2IX1 U2583 ( .B(res_not_wire[38]), .A(n3037), .Z(n3365) );
  CNR2IX1 U2584 ( .B(res_not_wire[36]), .A(n3033), .Z(n3682) );
  CNR2IX1 U2585 ( .B(n2965), .A(n3037), .Z(n3684) );
  CNR2IX1 U2586 ( .B(res_not_wire[32]), .A(n3037), .Z(n3686) );
  CND3XL U2587 ( .A(n1119), .B(n2141), .C(n56), .Z(n2250) );
  COND1XL U2588 ( .A(i[12]), .B(n3042), .C(n2202), .Z(n2204) );
  CENX1 U2589 ( .A(opera1[18]), .B(n2860), .Z(n3381) );
  CENX1 U2590 ( .A(opera1[19]), .B(n2860), .Z(n3388) );
  CNR3XL U2591 ( .A(n3699), .B(n56), .C(n2141), .Z(n2834) );
  COND11XL U2592 ( .A(n3042), .B(i[12]), .C(n2200), .D(n2201), .Z(n942) );
  COND11X1 U2593 ( .A(n3041), .B(i[14]), .C(n2145), .D(n2205), .Z(n940) );
  COND4CX1 U2594 ( .A(n3044), .B(n2152), .C(n2204), .D(i[14]), .Z(n2205) );
  COND11X1 U2595 ( .A(n3041), .B(i[27]), .C(n2100), .D(n2237), .Z(n927) );
  CND2X1 U2596 ( .A(i[27]), .B(n2238), .Z(n2237) );
  COND11X1 U2597 ( .A(n2230), .B(n2106), .C(n3042), .D(n2231), .Z(n930) );
  COND4CX1 U2598 ( .A(n3044), .B(n2106), .C(n2229), .D(i[24]), .Z(n2231) );
  COND1XL U2599 ( .A(n164), .B(n3037), .C(n2264), .Z(n918) );
  CANR2X1 U2600 ( .A(result[1]), .B(n3027), .C(n3021), .D(n2067), .Z(n2264) );
  COND1XL U2601 ( .A(n3034), .B(n2159), .C(n2272), .Z(n910) );
  CANR2X1 U2602 ( .A(result[9]), .B(n3027), .C(n3021), .D(n2063), .Z(n2272) );
  COND1XL U2603 ( .A(n3033), .B(n2138), .C(n2257), .Z(n920) );
  CANR2X1 U2604 ( .A(result[0]), .B(n3027), .C(n3021), .D(n3694), .Z(n2257) );
  COND1XL U2605 ( .A(n150), .B(n3038), .C(n2278), .Z(n904) );
  CANR2X1 U2606 ( .A(result[15]), .B(n3028), .C(n3022), .D(n2060), .Z(n2278)
         );
  COND1XL U2607 ( .A(n160), .B(n3037), .C(n2268), .Z(n914) );
  CANR2X1 U2608 ( .A(result[5]), .B(n3027), .C(n3021), .D(n2065), .Z(n2268) );
  COND1XL U2609 ( .A(n3035), .B(n2133), .C(n2279), .Z(n903) );
  CANR2X1 U2610 ( .A(result[16]), .B(n3028), .C(n3022), .D(n2075), .Z(n2279)
         );
  COND1XL U2611 ( .A(n162), .B(n3038), .C(n2266), .Z(n916) );
  CANR2X1 U2612 ( .A(result[3]), .B(n3027), .C(n3021), .D(n2066), .Z(n2266) );
  COND1XL U2613 ( .A(n154), .B(n3038), .C(n2274), .Z(n908) );
  CANR2X1 U2614 ( .A(result[11]), .B(n3027), .C(n3021), .D(n2062), .Z(n2274)
         );
  COND1XL U2615 ( .A(n3036), .B(n3698), .C(n2283), .Z(n899) );
  CANR2X1 U2616 ( .A(result[20]), .B(n3028), .C(n3022), .D(n2073), .Z(n2283)
         );
  COND1XL U2617 ( .A(n3035), .B(n2126), .C(n2285), .Z(n897) );
  CANR2X1 U2618 ( .A(result[22]), .B(n3028), .C(n3022), .D(n2072), .Z(n2285)
         );
  COND1XL U2619 ( .A(n3036), .B(n2124), .C(n2287), .Z(n895) );
  CANR2X1 U2620 ( .A(result[24]), .B(n3029), .C(n3023), .D(n2071), .Z(n2287)
         );
  COND1XL U2621 ( .A(n148), .B(n3038), .C(n2280), .Z(n902) );
  CANR2X1 U2622 ( .A(result[17]), .B(n3028), .C(n3022), .D(n2059), .Z(n2280)
         );
  COND1XL U2623 ( .A(n3034), .B(n2116), .C(n2297), .Z(n885) );
  COND1XL U2624 ( .A(n3036), .B(n3697), .C(n2289), .Z(n893) );
  CANR2X1 U2625 ( .A(result[26]), .B(n3029), .C(n3023), .D(n2070), .Z(n2289)
         );
  COND1XL U2626 ( .A(n3036), .B(n2110), .C(n2291), .Z(n891) );
  CANR2X1 U2627 ( .A(result[28]), .B(n3029), .C(n3023), .D(n2069), .Z(n2291)
         );
  COND1XL U2628 ( .A(n138), .B(n3039), .C(n2290), .Z(n892) );
  CANR2X1 U2629 ( .A(result[27]), .B(n3029), .C(n3023), .D(n2054), .Z(n2290)
         );
  COND1XL U2630 ( .A(n136), .B(n3039), .C(n2292), .Z(n890) );
  CANR2X1 U2631 ( .A(result[29]), .B(n3029), .C(n3023), .D(n2053), .Z(n2292)
         );
  COND1XL U2632 ( .A(n126), .B(n3039), .C(n2302), .Z(n880) );
  CANR2X1 U2633 ( .A(result[39]), .B(n3029), .C(n3023), .D(n2963), .Z(n2302)
         );
  COND1XL U2634 ( .A(n3035), .B(n2096), .C(n2303), .Z(n879) );
  CANR2X1 U2635 ( .A(result[40]), .B(n3030), .C(n3024), .D(n2955), .Z(n2303)
         );
  COND1XL U2636 ( .A(n3035), .B(n2095), .C(n2305), .Z(n877) );
  CANR2X1 U2637 ( .A(result[42]), .B(n3030), .C(n3024), .D(n2044), .Z(n2305)
         );
  COND1XL U2638 ( .A(n3035), .B(n2094), .C(n2309), .Z(n873) );
  CANR2X1 U2639 ( .A(result[46]), .B(n3030), .C(n3024), .D(n2040), .Z(n2309)
         );
  COND1XL U2640 ( .A(n124), .B(n3039), .C(n2304), .Z(n878) );
  CANR2X1 U2641 ( .A(result[41]), .B(n3030), .C(n3024), .D(n2045), .Z(n2304)
         );
  COND1XL U2642 ( .A(n3034), .B(n2091), .C(n2315), .Z(n867) );
  CANR2X1 U2643 ( .A(result[52]), .B(n3031), .C(n3025), .D(n2098), .Z(n2315)
         );
  COND1XL U2644 ( .A(n3034), .B(n3696), .C(n2313), .Z(n869) );
  CANR2X1 U2645 ( .A(result[50]), .B(n3030), .C(n3024), .D(n2038), .Z(n2313)
         );
  COND1XL U2646 ( .A(n114), .B(n3040), .C(n2314), .Z(n868) );
  CANR2X1 U2647 ( .A(result[51]), .B(n3030), .C(n3024), .D(n2097), .Z(n2314)
         );
  COND1XL U2648 ( .A(n112), .B(n3040), .C(n2316), .Z(n866) );
  CANR2X1 U2649 ( .A(result[53]), .B(n3031), .C(n3025), .D(n2036), .Z(n2316)
         );
  COND1XL U2650 ( .A(n3035), .B(n2088), .C(n2311), .Z(n871) );
  CANR2X1 U2651 ( .A(result[48]), .B(n3030), .C(n3024), .D(n2962), .Z(n2311)
         );
  COND1XL U2652 ( .A(n3033), .B(n2085), .C(n2324), .Z(n858) );
  CANR2X1 U2653 ( .A(result[61]), .B(n3031), .C(n3025), .D(n2032), .Z(n2324)
         );
  COND1XL U2654 ( .A(n3033), .B(n3674), .C(n2323), .Z(n859) );
  CANR2X1 U2655 ( .A(result[60]), .B(n3031), .C(n3025), .D(n2029), .Z(n2323)
         );
  COND1XL U2656 ( .A(n106), .B(n3037), .C(n2322), .Z(n860) );
  CANR2X1 U2657 ( .A(result[59]), .B(n3031), .C(n3025), .D(n2086), .Z(n2322)
         );
  COND1XL U2658 ( .A(n146), .B(n3038), .C(n2282), .Z(n900) );
  CANR2X1 U2659 ( .A(result[19]), .B(n3028), .C(n3022), .D(n2058), .Z(n2282)
         );
  COND1XL U2660 ( .A(n142), .B(n3038), .C(n2286), .Z(n896) );
  CANR2X1 U2661 ( .A(result[23]), .B(n3028), .C(n3022), .D(n2056), .Z(n2286)
         );
  COND1XL U2662 ( .A(n144), .B(n3038), .C(n2284), .Z(n898) );
  CANR2X1 U2663 ( .A(result[21]), .B(n3028), .C(n3022), .D(n2057), .Z(n2284)
         );
  COND1XL U2664 ( .A(n130), .B(n3039), .C(n2298), .Z(n884) );
  COND1XL U2665 ( .A(n140), .B(n3038), .C(n2288), .Z(n894) );
  CANR2X1 U2666 ( .A(result[25]), .B(n3029), .C(n3023), .D(n2055), .Z(n2288)
         );
  COND1XL U2667 ( .A(n134), .B(n3039), .C(n2294), .Z(n888) );
  CANR2X1 U2668 ( .A(result[31]), .B(n3029), .C(n3023), .D(n2051), .Z(n2294)
         );
  COND1XL U2669 ( .A(n120), .B(n3039), .C(n2308), .Z(n874) );
  CANR2X1 U2670 ( .A(result[45]), .B(n3030), .C(n3024), .D(n2113), .Z(n2308)
         );
  COND1XL U2671 ( .A(n122), .B(n3039), .C(n2306), .Z(n876) );
  CANR2X1 U2672 ( .A(result[43]), .B(n3030), .C(n3024), .D(n2046), .Z(n2306)
         );
  COND1XL U2673 ( .A(n116), .B(n3040), .C(n2312), .Z(n870) );
  CANR2X1 U2674 ( .A(result[49]), .B(n3030), .C(n3024), .D(n2961), .Z(n2312)
         );
  COND1XL U2675 ( .A(n110), .B(n3040), .C(n2318), .Z(n864) );
  CANR2X1 U2676 ( .A(result[55]), .B(n3031), .C(n3025), .D(n2092), .Z(n2318)
         );
  COND1XL U2677 ( .A(n118), .B(n3040), .C(n2310), .Z(n872) );
  CANR2X1 U2678 ( .A(result[47]), .B(n3030), .C(n3024), .D(n2112), .Z(n2310)
         );
  COND1XL U2679 ( .A(n3033), .B(n2031), .C(n2325), .Z(n857) );
  CANR2X1 U2680 ( .A(result[62]), .B(n3031), .C(n3025), .D(n3695), .Z(n2325)
         );
  COND1XL U2681 ( .A(n3034), .B(n3648), .C(n2320), .Z(n862) );
  CANR2X1 U2682 ( .A(result[57]), .B(n3031), .C(n3025), .D(n2033), .Z(n2320)
         );
  COND1XL U2683 ( .A(n3034), .B(n3693), .C(n2321), .Z(n861) );
  CANR2X1 U2684 ( .A(result[58]), .B(n3031), .C(n3025), .D(n2034), .Z(n2321)
         );
  COND1XL U2685 ( .A(n128), .B(n3039), .C(n2300), .Z(n882) );
  CANR2X1 U2686 ( .A(result[37]), .B(n3029), .C(n3023), .D(n2042), .Z(n2300)
         );
  COND1XL U2687 ( .A(n3035), .B(n3692), .C(n2307), .Z(n875) );
  CANR2X1 U2688 ( .A(result[44]), .B(n3030), .C(n3024), .D(n2115), .Z(n2307)
         );
  COND1XL U2689 ( .A(n3034), .B(n3702), .C(n2319), .Z(n863) );
  CANR2X1 U2690 ( .A(result[56]), .B(n3031), .C(n3025), .D(n2093), .Z(n2319)
         );
  COND1XL U2691 ( .A(n158), .B(n3038), .C(n2270), .Z(n912) );
  CANR2X1 U2692 ( .A(result[7]), .B(n3027), .C(n3021), .D(n2064), .Z(n2270) );
  COND1XL U2693 ( .A(n3033), .B(n2023), .C(n2269), .Z(n913) );
  CANR2X1 U2694 ( .A(result[6]), .B(n3027), .C(n3021), .D(n2052), .Z(n2269) );
  COND1XL U2695 ( .A(n2170), .B(n2156), .C(n2183), .Z(n950) );
  CND4XL U2696 ( .A(i[1]), .B(n3044), .C(n2156), .D(i[0]), .Z(n2183) );
  COND1XL U2697 ( .A(n2005), .B(n2152), .C(n2203), .Z(n941) );
  COND1XL U2698 ( .A(n3034), .B(n2147), .C(n2275), .Z(n907) );
  CANR2X1 U2699 ( .A(result[12]), .B(n3028), .C(n3022), .D(n2077), .Z(n2275)
         );
  COND4CX1 U2700 ( .A(n2232), .B(n2235), .C(n2121), .D(n2236), .Z(n928) );
  CND2X1 U2701 ( .A(n3044), .B(n2103), .Z(n2235) );
  COND4CX1 U2702 ( .A(n2242), .B(n2244), .C(n2104), .D(n2245), .Z(n924) );
  CND2X1 U2703 ( .A(n3044), .B(n2120), .Z(n2244) );
  CND4X1 U2704 ( .A(i[29]), .B(n3044), .C(n2104), .D(n3700), .Z(n2245) );
  COND1XL U2705 ( .A(n3036), .B(n2125), .C(n2281), .Z(n901) );
  CANR2X1 U2706 ( .A(result[18]), .B(n3028), .C(n3022), .D(n2074), .Z(n2281)
         );
  CND3XL U2707 ( .A(n2175), .B(n2174), .C(n2176), .Z(n953) );
  COND4CX1 U2708 ( .A(n3044), .B(n2155), .C(n2177), .D(i[5]), .Z(n2176) );
  CND2X1 U2709 ( .A(valid), .B(n3690), .Z(n2252) );
  CNR2IX1 U2710 ( .B(n960), .A(n3036), .Z(n3176) );
  CANR2X1 U2711 ( .A(result[13]), .B(n3028), .C(n3022), .D(n2061), .Z(n2276)
         );
  CNR2IX1 U2712 ( .B(res_not_wire[10]), .A(n3037), .Z(n3177) );
  CANR2X1 U2713 ( .A(result[10]), .B(n3027), .C(n3021), .D(n2078), .Z(n2273)
         );
  CNR2IXL U2714 ( .B(res_not_wire[2]), .A(n3037), .Z(n3178) );
  CANR2X1 U2715 ( .A(result[2]), .B(n3027), .C(n3021), .D(n2081), .Z(n2265) );
  CNR2IX1 U2716 ( .B(res_not_wire[8]), .A(n3036), .Z(n3212) );
  CANR2X1 U2717 ( .A(result[8]), .B(n3027), .C(n3021), .D(n2079), .Z(n2271) );
  CNR2IX1 U2718 ( .B(res_not_wire[14]), .A(n3036), .Z(n3213) );
  CANR2X1 U2719 ( .A(result[14]), .B(n3028), .C(n3022), .D(n2076), .Z(n2277)
         );
  CNR2IX1 U2720 ( .B(res_not_wire[4]), .A(n3037), .Z(n3687) );
  CANR2X1 U2721 ( .A(result[4]), .B(n3027), .C(n3021), .D(n2080), .Z(n2267) );
  CND2X1 U2722 ( .A(n2188), .B(n2189), .Z(n947) );
  COND4CX1 U2723 ( .A(n3044), .B(n2163), .C(n2187), .D(i[7]), .Z(n2188) );
  CND2X1 U2724 ( .A(n2193), .B(n2194), .Z(n945) );
  COND4CX1 U2725 ( .A(n3044), .B(n2143), .C(n2192), .D(i[9]), .Z(n2193) );
  CND2X1 U2726 ( .A(n2198), .B(n2199), .Z(n943) );
  COND4CX1 U2727 ( .A(n3044), .B(n2154), .C(n2197), .D(i[11]), .Z(n2198) );
  CND2X1 U2728 ( .A(n2210), .B(n2211), .Z(n938) );
  COND4CX1 U2729 ( .A(n3044), .B(n2129), .C(n2209), .D(i[16]), .Z(n2210) );
  CND2X1 U2730 ( .A(n2220), .B(n2221), .Z(n934) );
  COND4CX1 U2731 ( .A(n3044), .B(n2123), .C(n2219), .D(i[20]), .Z(n2220) );
  CND2X1 U2732 ( .A(n2215), .B(n2216), .Z(n936) );
  COND4CX1 U2733 ( .A(n3044), .B(n2119), .C(n2214), .D(i[18]), .Z(n2215) );
  CND2X1 U2734 ( .A(n2225), .B(n2226), .Z(n932) );
  COND4CX1 U2735 ( .A(n3044), .B(n2122), .C(n2224), .D(i[22]), .Z(n2225) );
  CND2X1 U2736 ( .A(n2239), .B(n2240), .Z(n926) );
  COND4CX1 U2737 ( .A(n3044), .B(n2102), .C(n2238), .D(i[28]), .Z(n2239) );
  CENX1 U2738 ( .A(n960), .B(n2988), .Z(n3118) );
  CEOX1 U2739 ( .A(opera2[17]), .B(n2002), .Z(n2744) );
  CENX1 U2740 ( .A(opera1[20]), .B(n2860), .Z(n3375) );
  CENX1 U2741 ( .A(opera1[21]), .B(n2860), .Z(n3373) );
  CENX1 U2742 ( .A(opera1[22]), .B(n2860), .Z(n3420) );
  CENX1 U2743 ( .A(opera1[24]), .B(n2860), .Z(n3430) );
  COND1XL U2744 ( .A(i[0]), .B(n3043), .C(n2178), .Z(n2182) );
  COND11XL U2745 ( .A(n3042), .B(i[8]), .C(n2190), .D(n2191), .Z(n946) );
  CND2X1 U2746 ( .A(i[8]), .B(n2192), .Z(n2191) );
  COND11XL U2747 ( .A(n3041), .B(i[6]), .C(n2185), .D(n2186), .Z(n948) );
  CND2X1 U2748 ( .A(i[6]), .B(n2187), .Z(n2186) );
  CND2XL U2749 ( .A(i[1]), .B(n2182), .Z(n2181) );
  COND11XL U2750 ( .A(n3041), .B(i[4]), .C(n2180), .D(n2184), .Z(n949) );
  CND2X1 U2751 ( .A(i[4]), .B(n2177), .Z(n2184) );
  COND11XL U2752 ( .A(n3042), .B(i[10]), .C(n2195), .D(n2196), .Z(n944) );
  CND2X1 U2753 ( .A(i[10]), .B(n2197), .Z(n2196) );
  COND11XL U2754 ( .A(n3041), .B(i[15]), .C(n2207), .D(n2208), .Z(n939) );
  CND2X1 U2755 ( .A(i[15]), .B(n2209), .Z(n2208) );
  COND11XL U2756 ( .A(n3041), .B(i[19]), .C(n2217), .D(n2218), .Z(n935) );
  CND2X1 U2757 ( .A(i[19]), .B(n2219), .Z(n2218) );
  COND11XL U2758 ( .A(n3041), .B(i[21]), .C(n2222), .D(n2223), .Z(n933) );
  CND2X1 U2759 ( .A(i[21]), .B(n2224), .Z(n2223) );
  COND11XL U2760 ( .A(n3041), .B(i[17]), .C(n2212), .D(n2213), .Z(n937) );
  CND2X1 U2761 ( .A(i[17]), .B(n2214), .Z(n2213) );
  COND11XL U2762 ( .A(n3041), .B(i[23]), .C(n2227), .D(n2228), .Z(n931) );
  CND2X1 U2763 ( .A(i[23]), .B(n2229), .Z(n2228) );
  COND2XL U2764 ( .A(n2162), .B(n2178), .C(i[0]), .D(n3041), .Z(n952) );
  CND3XL U2765 ( .A(res_not_wire[38]), .B(n3575), .C(n3226), .Z(n3306) );
  CND3XL U2766 ( .A(n53), .B(n2178), .C(n56), .Z(n2174) );
  COND1XL U2767 ( .A(n2140), .B(n3691), .C(n2164), .Z(n957) );
  CANR2X1 U2768 ( .A(n3690), .B(n2016), .C(nst[0]), .D(n2166), .Z(n2164) );
  COND1XL U2769 ( .A(n2250), .B(n2101), .C(n2251), .Z(n921) );
  CANR2X1 U2770 ( .A(n3690), .B(n2016), .C(nst[2]), .D(n2166), .Z(n2251) );
  CIVX2 U2771 ( .A(result[61]), .Z(n2032) );
  CENX1 U2772 ( .A(n3056), .B(res_not_wire[10]), .Z(n3128) );
  CENX1 U2773 ( .A(opera1[25]), .B(n2860), .Z(n3438) );
  CENX1 U2774 ( .A(opera1[26]), .B(n2860), .Z(n3473) );
  CENX1 U2775 ( .A(opera1[27]), .B(n2860), .Z(n3471) );
  CENX1 U2776 ( .A(opera1[28]), .B(n2860), .Z(n3484) );
  CENX1 U2777 ( .A(opera1[29]), .B(n2860), .Z(n3469) );
  CEOX1 U2778 ( .A(opera2[20]), .B(n2002), .Z(n2763) );
  CEOX1 U2779 ( .A(opera2[23]), .B(n2002), .Z(n2782) );
  COND1XL U2780 ( .A(n2016), .B(n2049), .C(n2249), .Z(n922) );
  CIVX2 U2781 ( .A(result[62]), .Z(n3695) );
  CENX1 U2782 ( .A(n162), .B(n3149), .Z(n3150) );
  CENX1 U2783 ( .A(n158), .B(n3137), .Z(n3138) );
  CENX1 U2784 ( .A(opera1[30]), .B(n2860), .Z(n3492) );
  CEOX1 U2785 ( .A(opera2[26]), .B(n2002), .Z(n2801) );
  CEOX1 U2786 ( .A(n2881), .B(n2860), .Z(n3179) );
  CNR2X1 U2787 ( .A(n2878), .B(nst[0]), .Z(n55) );
  CND2X1 U2788 ( .A(result[63]), .B(n3009), .Z(n3511) );
  CANR1XL U2789 ( .A(result[63]), .B(n3669), .C(n3459), .Z(n3500) );
  CANR2X1 U2790 ( .A(result[63]), .B(n3031), .C(n3025), .D(n3703), .Z(n2838)
         );
  CIVXL U2791 ( .A(n2241), .Z(n2100) );
  COND1XL U2792 ( .A(n2241), .B(n3042), .C(n2178), .Z(n2238) );
  CNIVXL U2793 ( .A(n3649), .Z(n2989) );
  CIVX3 U2794 ( .A(n3083), .Z(n3081) );
  CENX1 U2795 ( .A(opera1[4]), .B(opera1[31]), .Z(n3199) );
  CND2X1 U2796 ( .A(n3647), .B(n3646), .Z(n830) );
  CNR3XL U2797 ( .A(n3611), .B(n116), .C(n3696), .Z(n2983) );
  CIVX2 U2798 ( .A(n3158), .Z(n2984) );
  CND2X1 U2799 ( .A(n2720), .B(n2721), .Z(n811) );
  CIVX2 U2800 ( .A(n3117), .Z(n2985) );
  CIVX2 U2801 ( .A(n3649), .Z(n2986) );
  CANR2X1 U2802 ( .A(n2767), .B(n3688), .C(n2851), .D(n3092), .Z(n2766) );
  CENXL U2803 ( .A(n3504), .B(n3503), .Z(n3505) );
  COND2X1 U2804 ( .A(n3328), .B(n2113), .C(n3327), .D(n3326), .Z(n3346) );
  CNR2X1 U2805 ( .A(n3199), .B(n3198), .Z(n3200) );
  CNR2IXL U2806 ( .B(res_not_wire[18]), .A(n3105), .Z(n2990) );
  CNR2IX2 U2807 ( .B(res_not_wire[18]), .A(n3105), .Z(n2991) );
  CND2X1 U2808 ( .A(n3181), .B(n3180), .Z(n3189) );
  CNR2XL U2809 ( .A(n3067), .B(n2993), .Z(n2992) );
  CEOXL U2810 ( .A(n2674), .B(n2669), .Z(n2672) );
  CEOXL U2811 ( .A(n2655), .B(n2650), .Z(n2653) );
  CEOXL U2812 ( .A(n2788), .B(n2783), .Z(n2786) );
  CEOXL U2813 ( .A(n2807), .B(n2802), .Z(n2805) );
  CANR4CXL U2814 ( .A(n2795), .B(n2794), .C(n2801), .D(n2802), .Z(n2798) );
  CANR4CXL U2815 ( .A(n2776), .B(n2775), .C(n2782), .D(n2783), .Z(n2779) );
  CANR4CXL U2816 ( .A(n2662), .B(n2661), .C(n2668), .D(n2669), .Z(n2665) );
  CANR4CXL U2817 ( .A(n2642), .B(n2918), .C(n2649), .D(n2650), .Z(n2646) );
  CIVX2 U2818 ( .A(n3630), .Z(n2994) );
  CND2X1 U2819 ( .A(n3632), .B(n3631), .Z(n3639) );
  CNR2IXL U2820 ( .B(res_not_wire[52]), .A(n3409), .Z(n2995) );
  CNR2IX2 U2821 ( .B(res_not_wire[52]), .A(n3409), .Z(n3006) );
  CND2IX2 U2822 ( .B(n112), .A(n3006), .Z(n3630) );
  CAN2X1 U2823 ( .A(n3446), .B(res_not_wire[54]), .Z(n2997) );
  CANR4CXL U2824 ( .A(n2757), .B(n2756), .C(n2763), .D(n2764), .Z(n2760) );
  CIVX2 U2825 ( .A(n3056), .Z(n2999) );
  CEOXL U2826 ( .A(n3671), .B(n3670), .Z(n3672) );
  CENXL U2827 ( .A(n3418), .B(n3416), .Z(n3396) );
  CNR2IXL U2828 ( .B(n2948), .A(n3260), .Z(n3264) );
  CENX1 U2829 ( .A(opera1[3]), .B(opera1[31]), .Z(n3198) );
  CENX1 U2830 ( .A(opera1[2]), .B(opera1[31]), .Z(n3196) );
  CND2IX2 U2831 ( .B(n3002), .A(n3052), .Z(n3140) );
  COR4X1 U2832 ( .A(n3308), .B(n3307), .C(n3306), .D(n124), .Z(n3004) );
  COND2X1 U2833 ( .A(n2137), .B(n2167), .C(n3179), .D(n2004), .Z(n956) );
  CENX1 U2834 ( .A(result[63]), .B(n3497), .Z(n3498) );
  COND1XL U2835 ( .A(n3525), .B(n3253), .C(n3255), .Z(n3563) );
  CND2XL U2836 ( .A(result[36]), .B(n3195), .Z(n3255) );
  CENX1 U2837 ( .A(result[36]), .B(n3195), .Z(n3253) );
  CND2IXL U2838 ( .B(n3141), .A(n3140), .Z(n3142) );
  CND2IXL U2839 ( .B(n2848), .A(n3510), .Z(n3501) );
  CND2X1 U2840 ( .A(res_not_wire[14]), .B(n960), .Z(n3005) );
  CENX1 U2841 ( .A(n3510), .B(n2050), .Z(n3512) );
  CND3XL U2842 ( .A(n3677), .B(n3676), .C(n2849), .Z(n3678) );
  CND2IXL U2843 ( .B(n3122), .A(n3121), .Z(n3123) );
  CND3XL U2844 ( .A(n2851), .B(n3651), .C(n3650), .Z(n3658) );
  CND2IXL U2845 ( .B(n3354), .A(n3353), .Z(n3355) );
  COND1XL U2846 ( .A(n2989), .B(n3702), .C(n3648), .Z(n3650) );
  CNR2IXL U2847 ( .B(n3083), .A(n2848), .Z(n3089) );
  COND1XL U2848 ( .A(n3131), .B(n158), .C(n3130), .Z(n3132) );
  COND1XL U2849 ( .A(n2987), .B(n164), .C(n3151), .Z(n3152) );
  CND2IXL U2850 ( .B(res_not_wire[58]), .A(n3651), .Z(n3644) );
  CND2IXL U2851 ( .B(n3103), .A(n3102), .Z(n3104) );
  CND2IXL U2852 ( .B(res_not_wire[48]), .A(n3310), .Z(n3340) );
  CNR2IXL U2853 ( .B(n3075), .A(n2850), .Z(n3077) );
  CANR1XL U2854 ( .A(n1053), .B(n3659), .C(res_not_wire[62]), .Z(n3502) );
  COND3XL U2855 ( .A(n2995), .B(n2871), .C(n2851), .D(n2996), .Z(n3629) );
  CANR11XL U2856 ( .A(n3116), .B(n3115), .C(n2849), .D(n2864), .Z(n2721) );
  CND2IXL U2857 ( .B(res_not_wire[54]), .A(n2996), .Z(n3631) );
  CND2IXL U2858 ( .B(n3085), .A(n3084), .Z(n3088) );
  CND3XL U2859 ( .A(n2851), .B(n3153), .C(n3152), .Z(n3156) );
  CND2IXL U2860 ( .B(res_not_wire[30]), .A(n3067), .Z(n3065) );
  CNR2IXL U2861 ( .B(n136), .A(n3001), .Z(n3068) );
  CNR2IXL U2862 ( .B(n3067), .A(n2852), .Z(n3070) );
  CNR3XL U2863 ( .A(n2857), .B(n1061), .C(n2250), .Z(n2258) );
  CND2IXL U2864 ( .B(n2850), .A(n3524), .Z(n3531) );
  CNR2IXL U2865 ( .B(n2849), .A(n3352), .Z(n3356) );
  COND3X1 U2866 ( .A(n3509), .B(n2850), .C(n3508), .D(n3507), .Z(n829) );
  CND3XL U2867 ( .A(n2847), .B(n3124), .C(n3123), .Z(n3127) );
  CND3XL U2868 ( .A(n2849), .B(n3143), .C(n3142), .Z(n3146) );
  CND2IXL U2869 ( .B(res_not_wire[36]), .A(n3524), .Z(n3207) );
  CND2IXL U2870 ( .B(n146), .A(n2990), .Z(n3093) );
  CNR2IXL U2871 ( .B(n2849), .A(n2998), .Z(n3632) );
  CNR2IXL U2872 ( .B(n2851), .A(n3000), .Z(n3181) );
  CNR2IXL U2873 ( .B(n2847), .A(n2983), .Z(n3603) );
  CANR1XL U2874 ( .A(res_not_wire[34]), .B(n3000), .C(n3523), .Z(n3532) );
  CANR11XL U2875 ( .A(n2849), .B(n3611), .C(n3340), .D(n3339), .Z(n3343) );
  CANR11XL U2876 ( .A(n2851), .B(n3222), .C(n3221), .D(n3220), .Z(n3223) );
  CND2IXL U2877 ( .B(n2965), .A(n3222), .Z(n3180) );
  COND1XL U2878 ( .A(n3611), .B(n116), .C(n3696), .Z(n3602) );
  CND3XL U2879 ( .A(n2849), .B(n3105), .C(n3104), .Z(n3108) );
  COND1XL U2880 ( .A(n3675), .B(n106), .C(n3674), .Z(n3676) );
  CND3XL U2881 ( .A(n2851), .B(n3133), .C(n3132), .Z(n3136) );
  CND3XL U2882 ( .A(n2847), .B(n3095), .C(n3094), .Z(n3098) );
  COND1XL U2883 ( .A(n2988), .B(n3114), .C(n3113), .Z(n3115) );
  CND2IXL U2884 ( .B(n134), .A(n2992), .Z(n3219) );
  CNR2XL U2885 ( .A(n2992), .B(n2848), .Z(n3066) );
  COND1XL U2886 ( .A(n3079), .B(n140), .C(n3697), .Z(n3076) );
  CND2IX2 U2887 ( .B(n3050), .A(n3049), .Z(n3668) );
  CND2X4 U2888 ( .A(result[0]), .B(n3689), .Z(n3673) );
  CIVXL U2889 ( .A(n3012), .Z(n3009) );
  CIVXL U2890 ( .A(n2857), .Z(n3033) );
  CIVXL U2891 ( .A(n2857), .Z(n3035) );
  CIVXL U2892 ( .A(n2857), .Z(n3036) );
  CIVXL U2893 ( .A(n2857), .Z(n3040) );
  CIVXL U2894 ( .A(n3043), .Z(n3044) );
  CAN2X1 U2895 ( .A(n53), .B(n56), .Z(n3045) );
  CND2IX1 U2896 ( .B(n1119), .A(n3045), .Z(n3064) );
  CIVX2 U2897 ( .A(n3064), .Z(n3690) );
  CIVX2 U2898 ( .A(n2883), .Z(n3691) );
  CIVX2 U2899 ( .A(n2250), .Z(n3701) );
  CIVX2 U2900 ( .A(n3048), .Z(n2169) );
  CIVX2 U2901 ( .A(result[63]), .Z(n3703) );
  CIVX2 U2902 ( .A(n1056), .Z(n2050) );
  CND2IX1 U2903 ( .B(n2247), .A(n3048), .Z(n3049) );
  CND2IX1 U2904 ( .B(n2250), .A(n3020), .Z(n3051) );
  CIVX2 U2905 ( .A(n3051), .Z(n3689) );
  CND2IX1 U2906 ( .B(n2140), .A(n3019), .Z(n3086) );
  CIVX2 U2907 ( .A(n136), .Z(n3063) );
  CIVX2 U2908 ( .A(n140), .Z(n3078) );
  CIVX2 U2909 ( .A(res_not_wire[26]), .Z(n3697) );
  CIVX2 U2910 ( .A(n142), .Z(n3085) );
  CIVX2 U2911 ( .A(n144), .Z(n3091) );
  CIVX2 U2912 ( .A(n148), .Z(n3103) );
  CIVX2 U2913 ( .A(n154), .Z(n3122) );
  CIVX2 U2914 ( .A(n164), .Z(n3157) );
  CIVX2 U2915 ( .A(n3153), .Z(n3149) );
  CIVX2 U2916 ( .A(n3147), .Z(n3052) );
  CIVX2 U2917 ( .A(n3140), .Z(n3053) );
  CIVX2 U2918 ( .A(n3143), .Z(n3054) );
  CND2X2 U2919 ( .A(n3054), .B(res_not_wire[6]), .Z(n3131) );
  CIVX2 U2920 ( .A(n3133), .Z(n3055) );
  CND2X2 U2921 ( .A(n962), .B(n3055), .Z(n3056) );
  CND2X2 U2922 ( .A(n2999), .B(res_not_wire[10]), .Z(n3121) );
  CIVX2 U2923 ( .A(n3121), .Z(n3057) );
  CND2X2 U2924 ( .A(res_not_wire[12]), .B(n3119), .Z(n3117) );
  CND2X2 U2925 ( .A(n2867), .B(n3111), .Z(n3109) );
  CIVX2 U2926 ( .A(n3109), .Z(n3058) );
  CIVX2 U2927 ( .A(n3102), .Z(n3059) );
  CND2X2 U2928 ( .A(n3103), .B(n3059), .Z(n3105) );
  CND2X2 U2929 ( .A(n2925), .B(res_not_wire[22]), .Z(n3084) );
  CIVX2 U2930 ( .A(n3084), .Z(n3060) );
  CND2X2 U2931 ( .A(n3085), .B(n3060), .Z(n3083) );
  CND2X2 U2932 ( .A(res_not_wire[24]), .B(n3081), .Z(n3079) );
  CIVX2 U2933 ( .A(n3079), .Z(n3061) );
  CANR2X1 U2934 ( .A(n2824), .B(n3688), .C(n3066), .D(n3065), .Z(n2823) );
  CIVX2 U2935 ( .A(n3068), .Z(n3069) );
  CANR2X1 U2936 ( .A(n2817), .B(n3688), .C(n3070), .D(n3069), .Z(n2816) );
  CANR2X1 U2937 ( .A(n2810), .B(n3688), .C(n2849), .D(n3072), .Z(n2809) );
  CANR2X1 U2938 ( .A(n2805), .B(n3688), .C(n2849), .D(n3074), .Z(n2804) );
  CANR2X1 U2939 ( .A(n2798), .B(n3688), .C(n3077), .D(n3076), .Z(n2797) );
  CIVX2 U2940 ( .A(res_not_wire[22]), .Z(n2126) );
  CND2IX1 U2941 ( .B(res_not_wire[20]), .A(n3093), .Z(n3094) );
  CIVX2 U2942 ( .A(n2760), .Z(n3096) );
  CND2IX1 U2943 ( .B(n3096), .A(n3688), .Z(n3097) );
  CAN2X1 U2944 ( .A(n3098), .B(n3097), .Z(n2759) );
  CIVX2 U2945 ( .A(n2125), .Z(n3100) );
  CIVX2 U2946 ( .A(n2741), .Z(n3106) );
  CND2IX1 U2947 ( .B(n3106), .A(n3688), .Z(n3107) );
  CAN2X1 U2948 ( .A(n3108), .B(n3107), .Z(n2740) );
  CIVX2 U2949 ( .A(n960), .Z(n3114) );
  CIVX2 U2950 ( .A(res_not_wire[14]), .Z(n3113) );
  CIVX2 U2951 ( .A(n2703), .Z(n3125) );
  CND2IX1 U2952 ( .B(n3125), .A(n3688), .Z(n3126) );
  CAN2X1 U2953 ( .A(n3127), .B(n3126), .Z(n2702) );
  CIVX2 U2954 ( .A(res_not_wire[8]), .Z(n3130) );
  CIVX2 U2955 ( .A(n2684), .Z(n3134) );
  CND2IX1 U2956 ( .B(n3134), .A(n3688), .Z(n3135) );
  CAN2X1 U2957 ( .A(n3136), .B(n3135), .Z(n2683) );
  CIVX2 U2958 ( .A(n2665), .Z(n3144) );
  CND2IX1 U2959 ( .B(n3144), .A(n3688), .Z(n3145) );
  CAN2X1 U2960 ( .A(n3146), .B(n3145), .Z(n2664) );
  CIVX2 U2961 ( .A(res_not_wire[2]), .Z(n3151) );
  CIVX2 U2962 ( .A(n2646), .Z(n3154) );
  CND2IX1 U2963 ( .B(n3154), .A(n3688), .Z(n3155) );
  CAN2X1 U2964 ( .A(n3156), .B(n3155), .Z(n2645) );
  CIVX2 U2965 ( .A(res_not_wire[34]), .Z(n2116) );
  CENX1 U2966 ( .A(opera1[31]), .B(opera1[1]), .Z(n3162) );
  CND3X2 U2967 ( .A(c_inop1), .B(n2922), .C(n2956), .Z(n3165) );
  CIVX2 U2968 ( .A(n3165), .Z(n3202) );
  CIVX2 U2969 ( .A(n3196), .Z(n3160) );
  CIVX2 U2970 ( .A(n3168), .Z(n3183) );
  CIVX2 U2971 ( .A(n3514), .Z(n3513) );
  CND2X2 U2972 ( .A(result[32]), .B(n3513), .Z(n3214) );
  CIVX2 U2973 ( .A(n3214), .Z(n3167) );
  CND2IX1 U2974 ( .B(result[33]), .A(n3215), .Z(n3166) );
  CIVX2 U2975 ( .A(n3182), .Z(n3170) );
  CND2IX1 U2976 ( .B(result[34]), .A(n3168), .Z(n3169) );
  COND4CX1 U2977 ( .A(result[34]), .B(n3183), .C(n3170), .D(n3169), .Z(n3192)
         );
  CIVX2 U2978 ( .A(n3192), .Z(n3173) );
  CENX1 U2979 ( .A(n3173), .B(n3193), .Z(n3174) );
  CANR2X1 U2980 ( .A(n2847), .B(n3175), .C(n3642), .D(n3174), .Z(n2348) );
  CIVX2 U2981 ( .A(n1053), .Z(n2085) );
  CIVX2 U2982 ( .A(result[60]), .Z(n2029) );
  CIVX2 U2983 ( .A(result[59]), .Z(n2086) );
  CIVX2 U2984 ( .A(result[58]), .Z(n2034) );
  CIVX2 U2985 ( .A(res_not_wire[58]), .Z(n3693) );
  CIVX2 U2986 ( .A(result[57]), .Z(n2033) );
  CIVX2 U2987 ( .A(result[56]), .Z(n2093) );
  CIVX2 U2988 ( .A(res_not_wire[56]), .Z(n3702) );
  CIVX2 U2989 ( .A(result[55]), .Z(n2092) );
  CIVX2 U2990 ( .A(result[54]), .Z(n2035) );
  CIVX2 U2991 ( .A(result[53]), .Z(n2036) );
  CIVX2 U2992 ( .A(result[52]), .Z(n2098) );
  CIVX2 U2993 ( .A(res_not_wire[52]), .Z(n2091) );
  CIVX2 U2994 ( .A(result[51]), .Z(n2097) );
  CIVX2 U2995 ( .A(result[50]), .Z(n2038) );
  CIVX2 U2996 ( .A(res_not_wire[50]), .Z(n3696) );
  CIVX2 U2997 ( .A(result[47]), .Z(n2112) );
  CIVX2 U2998 ( .A(result[46]), .Z(n2040) );
  CIVX2 U2999 ( .A(res_not_wire[46]), .Z(n2094) );
  CIVX2 U3000 ( .A(result[45]), .Z(n2113) );
  CIVX2 U3001 ( .A(result[44]), .Z(n2115) );
  CIVX2 U3002 ( .A(res_not_wire[44]), .Z(n3692) );
  CIVX2 U3003 ( .A(result[43]), .Z(n2046) );
  CIVX2 U3004 ( .A(result[42]), .Z(n2044) );
  CIVX2 U3005 ( .A(res_not_wire[40]), .Z(n2096) );
  CIVX2 U3006 ( .A(res_not_wire[28]), .Z(n2110) );
  CIVX2 U3007 ( .A(res_not_wire[20]), .Z(n3698) );
  CIVX2 U3008 ( .A(res_not_wire[16]), .Z(n2133) );
  CIVX2 U3009 ( .A(n2246), .Z(n3700) );
  CND2IX1 U3010 ( .B(n3176), .A(n2276), .Z(n906) );
  CND2IX1 U3011 ( .B(n3177), .A(n2273), .Z(n909) );
  CND2IX1 U3012 ( .B(n3178), .A(n2265), .Z(n917) );
  CEO3X1 U3013 ( .A(n2047), .B(n3183), .C(n3182), .Z(n3184) );
  CIVX2 U3014 ( .A(n2047), .Z(n3186) );
  CIVX2 U3015 ( .A(n130), .Z(n3523) );
  CIVX2 U3016 ( .A(n3204), .Z(n3203) );
  CND2X2 U3017 ( .A(result[37]), .B(n3203), .Z(n3562) );
  CND2IX1 U3018 ( .B(result[37]), .A(n3204), .Z(n3205) );
  CND2X2 U3019 ( .A(n3562), .B(n3205), .Z(n3564) );
  CENX1 U3020 ( .A(n3563), .B(n3564), .Z(n3206) );
  CND2IX1 U3021 ( .B(n3212), .A(n2271), .Z(n911) );
  CND2IX1 U3022 ( .B(n3213), .A(n2277), .Z(n905) );
  CND2IX1 U3023 ( .B(n2920), .A(n3669), .Z(n3225) );
  CENX1 U3024 ( .A(result[33]), .B(n3215), .Z(n3216) );
  CMXI2X1 U3025 ( .A0(n3218), .A1(n3217), .S(n3216), .Z(n3224) );
  CND2IX1 U3026 ( .B(res_not_wire[32]), .A(n3219), .Z(n3221) );
  CIVX2 U3027 ( .A(n128), .Z(n3575) );
  CENX1 U3028 ( .A(n3541), .B(n2096), .Z(n3269) );
  CIVX2 U3029 ( .A(n3236), .Z(n3228) );
  CIVX2 U3030 ( .A(n3235), .Z(n3227) );
  CND2X2 U3031 ( .A(n3228), .B(n3227), .Z(n3240) );
  CIVX2 U3032 ( .A(n3240), .Z(n3230) );
  CIVX2 U3033 ( .A(n3239), .Z(n3229) );
  CIVX2 U3034 ( .A(n3242), .Z(n3232) );
  CIVX2 U3035 ( .A(n3233), .Z(n3231) );
  CND2X2 U3036 ( .A(n3232), .B(n3231), .Z(n3248) );
  CIVX2 U3037 ( .A(n3256), .Z(n3586) );
  CIVX2 U3038 ( .A(n3248), .Z(n3246) );
  CIVX2 U3039 ( .A(n3247), .Z(n3245) );
  CIVX2 U3040 ( .A(n3251), .Z(n3250) );
  CND2IX1 U3041 ( .B(result[41]), .A(n3251), .Z(n3252) );
  CIVX2 U3042 ( .A(n3253), .Z(n3526) );
  COND2X2 U3043 ( .A(n3255), .B(n3564), .C(n3254), .D(n3525), .Z(n3260) );
  CIVX2 U3044 ( .A(n3260), .Z(n3257) );
  CND2X1 U3045 ( .A(n3259), .B(n3258), .Z(n3278) );
  COND3X1 U3046 ( .A(n3269), .B(n2850), .C(n3268), .D(n3267), .Z(n848) );
  CIVX2 U3047 ( .A(n122), .Z(n3533) );
  CIVX2 U3048 ( .A(n3306), .Z(n3270) );
  CIVX2 U3049 ( .A(n124), .Z(n3542) );
  CND2IX1 U3050 ( .B(n2850), .A(n3344), .Z(n3304) );
  CIVX2 U3051 ( .A(n3280), .Z(n3272) );
  CIVX2 U3052 ( .A(n3279), .Z(n3271) );
  CIVX2 U3053 ( .A(n3282), .Z(n3274) );
  CIVX2 U3054 ( .A(n3275), .Z(n3273) );
  CIVX2 U3055 ( .A(n3544), .Z(n3285) );
  CIVX2 U3056 ( .A(n3290), .Z(n3288) );
  CIVX2 U3057 ( .A(n3289), .Z(n3287) );
  CIVX2 U3058 ( .A(n3534), .Z(n3294) );
  CIVX2 U3059 ( .A(n3298), .Z(n3296) );
  CIVX2 U3060 ( .A(n3297), .Z(n3295) );
  COND3X1 U3061 ( .A(n3305), .B(n3304), .C(n3303), .D(n3302), .Z(n844) );
  CIVX2 U3062 ( .A(n118), .Z(n3354) );
  CND4X1 U3063 ( .A(n2870), .B(res_not_wire[36]), .C(n3533), .D(
        res_not_wire[44]), .Z(n3308) );
  CND2X2 U3064 ( .A(res_not_wire[46]), .B(n3003), .Z(n3353) );
  CIVX2 U3065 ( .A(n3353), .Z(n3309) );
  CIVX2 U3066 ( .A(n3310), .Z(n3352) );
  CND2X2 U3067 ( .A(res_not_wire[48]), .B(n3352), .Z(n3611) );
  CIVX2 U3068 ( .A(n3323), .Z(n3312) );
  CIVX2 U3069 ( .A(n3322), .Z(n3311) );
  CIVX2 U3070 ( .A(n3325), .Z(n3314) );
  CIVX2 U3071 ( .A(n3319), .Z(n3313) );
  CIVX2 U3072 ( .A(n3321), .Z(n3316) );
  CIVX2 U3073 ( .A(n3317), .Z(n3315) );
  CIVX2 U3074 ( .A(n3345), .Z(n3331) );
  CANR1X2 U3075 ( .A(n3331), .B(n3346), .C(n3330), .Z(n3596) );
  CIVX2 U3076 ( .A(n3337), .Z(n3335) );
  CIVX2 U3077 ( .A(n3336), .Z(n3334) );
  CENX1 U3078 ( .A(n120), .B(n3344), .Z(n3351) );
  CMXI2X1 U3079 ( .A0(n3026), .A1(n3032), .S(result[38]), .Z(n3364) );
  CND2IX1 U3080 ( .B(n3365), .A(n3364), .Z(n881) );
  CIVX2 U3081 ( .A(n114), .Z(n3401) );
  CIVX2 U3082 ( .A(n3382), .Z(n3367) );
  CIVX2 U3083 ( .A(n3381), .Z(n3366) );
  CIVX2 U3084 ( .A(n3388), .Z(n3368) );
  CIVX2 U3085 ( .A(n3391), .Z(n3370) );
  CIVX2 U3086 ( .A(n3375), .Z(n3369) );
  CIVX2 U3087 ( .A(n3377), .Z(n3372) );
  CIVX2 U3088 ( .A(n3373), .Z(n3371) );
  CIVX2 U3089 ( .A(n3384), .Z(n3385) );
  CNR2X2 U3090 ( .A(n3394), .B(n3393), .Z(n3403) );
  COND2X2 U3091 ( .A(n3395), .B(n2098), .C(n3403), .D(n3402), .Z(n3416) );
  COND3X1 U3092 ( .A(n3400), .B(n2850), .C(n3399), .D(n3398), .Z(n836) );
  CIVX2 U3093 ( .A(n110), .Z(n3446) );
  CND2X2 U3094 ( .A(n2994), .B(n2997), .Z(n3649) );
  CIVX2 U3095 ( .A(n3421), .Z(n3411) );
  CIVX2 U3096 ( .A(n3420), .Z(n3410) );
  CIVX2 U3097 ( .A(n3423), .Z(n3413) );
  CIVX2 U3098 ( .A(n3414), .Z(n3412) );
  CIVX2 U3099 ( .A(n3416), .Z(n3417) );
  CIVX2 U3100 ( .A(n3623), .Z(n3426) );
  CANR1X2 U3101 ( .A(n3624), .B(n3426), .C(n3425), .Z(n3634) );
  COND2X2 U3102 ( .A(n3427), .B(n2092), .C(n3634), .D(n3633), .Z(n3448) );
  CIVX2 U3103 ( .A(n3431), .Z(n3429) );
  CIVX2 U3104 ( .A(n3430), .Z(n3428) );
  CANR1X2 U3105 ( .A(n3448), .B(n3435), .C(n3434), .Z(n3477) );
  CIVX2 U3106 ( .A(n3439), .Z(n3437) );
  CIVX2 U3107 ( .A(n3438), .Z(n3436) );
  COND3X1 U3108 ( .A(n3445), .B(n2852), .C(n3444), .D(n3443), .Z(n832) );
  CIVX2 U3109 ( .A(res_not_wire[60]), .Z(n3674) );
  CAN2X1 U3110 ( .A(n1093), .B(res_not_wire[56]), .Z(n3454) );
  CIVX2 U3111 ( .A(n3651), .Z(n3455) );
  CND2X2 U3112 ( .A(n3455), .B(res_not_wire[58]), .Z(n3675) );
  CIVX2 U3113 ( .A(n3675), .Z(n3456) );
  CND2X2 U3114 ( .A(n3456), .B(n3457), .Z(n3677) );
  CAN2X1 U3115 ( .A(res_not_wire[62]), .B(n1053), .Z(n3458) );
  CND2X2 U3116 ( .A(n3659), .B(n3458), .Z(n3510) );
  CIVX2 U3117 ( .A(n3492), .Z(n3460) );
  CIVX2 U3118 ( .A(n3474), .Z(n3462) );
  CIVX2 U3119 ( .A(n3473), .Z(n3461) );
  CIVX2 U3120 ( .A(n3476), .Z(n3464) );
  CIVX2 U3121 ( .A(n3471), .Z(n3463) );
  CIVX2 U3122 ( .A(n3485), .Z(n3466) );
  CIVX2 U3123 ( .A(n3484), .Z(n3465) );
  CIVX2 U3124 ( .A(n3487), .Z(n3468) );
  CIVX2 U3125 ( .A(n3469), .Z(n3467) );
  CIVX2 U3126 ( .A(n3660), .Z(n3496) );
  CIVX2 U3127 ( .A(n3652), .Z(n3482) );
  COND2X2 U3128 ( .A(n3483), .B(n2086), .C(n3641), .D(n3640), .Z(n3504) );
  CIVX2 U3129 ( .A(n3503), .Z(n3490) );
  CANR1X2 U3130 ( .A(n3504), .B(n3490), .C(n3489), .Z(n3670) );
  COND2X2 U3131 ( .A(n3491), .B(n2032), .C(n3670), .D(n3671), .Z(n3661) );
  CND2IX1 U3132 ( .B(n3673), .A(n3505), .Z(n3508) );
  CMXI2X1 U3133 ( .A0(n3517), .A1(n3516), .S(result[32]), .Z(n3518) );
  CND2IX1 U3134 ( .B(n3519), .A(n3518), .Z(n3522) );
  CANR2X1 U3135 ( .A(n2829), .B(n3688), .C(n2847), .D(n3520), .Z(n3521) );
  CENX1 U3136 ( .A(n3526), .B(n3525), .Z(n3527) );
  COND3X1 U3137 ( .A(n3532), .B(n3531), .C(n3530), .D(n3529), .Z(n853) );
  CENX1 U3138 ( .A(n2954), .B(n3533), .Z(n3540) );
  CENX1 U3139 ( .A(n3545), .B(n3544), .Z(n3546) );
  CND2IX1 U3140 ( .B(n2852), .A(n3583), .Z(n3573) );
  CIVX2 U3141 ( .A(n3576), .Z(n3567) );
  CND2IX1 U3142 ( .B(n3564), .A(n3563), .Z(n3584) );
  CIVX2 U3143 ( .A(n3565), .Z(n3566) );
  COND3X1 U3144 ( .A(n3574), .B(n3573), .C(n3572), .D(n3571), .Z(n850) );
  CENX1 U3145 ( .A(n2952), .B(n3575), .Z(n3582) );
  CENX1 U3146 ( .A(n3577), .B(n3576), .Z(n3578) );
  CENX1 U3147 ( .A(n126), .B(n3583), .Z(n3594) );
  CND2IX1 U3148 ( .B(n3585), .A(n3584), .Z(n3587) );
  COND3X1 U3149 ( .A(n3601), .B(n2848), .C(n3600), .D(n3599), .Z(n842) );
  CIVX2 U3150 ( .A(n3613), .Z(n3617) );
  CIVX2 U3151 ( .A(n3614), .Z(n3615) );
  CIVX2 U3152 ( .A(n1093), .Z(n3648) );
  CND2IX1 U3153 ( .B(n3673), .A(n3654), .Z(n3657) );
  CENX1 U3154 ( .A(n3661), .B(n3660), .Z(n3662) );
  CND2IX1 U3155 ( .B(n3673), .A(n3662), .Z(n3665) );
  COND3X1 U3156 ( .A(n3667), .B(n2848), .C(n3665), .D(n3664), .Z(n827) );
  CND2IX1 U3157 ( .B(n3673), .A(n3672), .Z(n3679) );
  CMXI2X1 U3158 ( .A0(n3026), .A1(n3032), .S(result[36]), .Z(n3681) );
  CND2IX1 U3159 ( .B(n3682), .A(n3681), .Z(n883) );
  CND2IX1 U3160 ( .B(n3684), .A(n3683), .Z(n886) );
  CND2IX1 U3161 ( .B(n3686), .A(n3685), .Z(n887) );
  CND2IX1 U3162 ( .B(n3687), .A(n2267), .Z(n915) );
endmodule



module multiplier ( result, valid, opera1, opera2, muordi, clock, reset, start
 );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input muordi, clock, reset, start;
  output valid;
  wire   opera2_63, N34, n52, n53, n55, n56, n106, n110, n112, n114, n116,
         n118, n120, n122, n124, n126, n128, n130, n134, n136, n138, n140,
         n142, n144, n146, n148, n150, n154, n158, n160, n162, n164, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n957, n960, n962,
         n1053, n1056, n1061, n1093, n1119, n2001, n2003, n2005, n2007, n2008,
         n2015, n2016, n2023, n2029, n2031, n2032, n2033, n2034, n2035, n2036,
         n2038, n2040, n2042, n2044, n2045, n2046, n2047, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2085, n2086, n2088, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2110,
         n2112, n2113, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2129, n2130, n2133, n2137, n2138, n2140,
         n2141, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2159, n2162, n2163, n2164,
         n2166, n2167, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2297, n2298, n2300, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2330, n2347, n2348, n2630, n2631, n2633, n2634, n2635, n2637, n2638,
         n2639, n2642, n2643, n2644, n2646, n2649, n2650, n2651, n2652, n2653,
         n2655, n2656, n2657, n2658, n2661, n2662, n2663, n2665, n2668, n2669,
         n2670, n2671, n2672, n2674, n2675, n2676, n2677, n2680, n2681, n2682,
         n2684, n2687, n2688, n2689, n2690, n2691, n2693, n2694, n2695, n2696,
         n2699, n2700, n2701, n2703, n2706, n2707, n2708, n2709, n2710, n2712,
         n2713, n2714, n2715, n2718, n2719, n2720, n2721, n2722, n2725, n2726,
         n2727, n2728, n2729, n2731, n2732, n2733, n2734, n2737, n2738, n2739,
         n2741, n2744, n2745, n2746, n2747, n2748, n2750, n2751, n2752, n2753,
         n2756, n2757, n2758, n2760, n2763, n2764, n2766, n2767, n2769, n2770,
         n2771, n2772, n2775, n2776, n2777, n2778, n2779, n2782, n2783, n2785,
         n2786, n2788, n2789, n2790, n2791, n2794, n2795, n2796, n2797, n2798,
         n2801, n2802, n2803, n2804, n2805, n2807, n2808, n2809, n2810, n2813,
         n2814, n2815, n2816, n2817, n2820, n2821, n2823, n2824, n2826, n2829,
         n2833, n2834, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2866, n2867, n2868, n2869, n2870, n2871, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588;
  wire   [63:0] res_not_wire;
  wire   [2:0] nst;
  wire   [31:0] i;
  tri   c_inop1;
  tri   c_inop2;
  tri   c_inres;
  assign opera2_63 = opera2[63];

  CTSX2 A4 ( .A(1'b0), .E(n2866), .Z(c_inop2) );
  CTSX2 A3 ( .A(1'b1), .E(opera2_63), .Z(c_inop2) );
  CTSX2 A6 ( .A(1'b0), .E(n2137), .Z(c_inres) );
  CTSX2 A5 ( .A(1'b1), .E(n1061), .Z(c_inres) );
  CIVX2 U1667 ( .A(n2821), .Z(n2001) );
  CIVX2 U1671 ( .A(n2204), .Z(n2005) );
  CIVX2 U1673 ( .A(n2178), .Z(n2007) );
  CIVX2 U1674 ( .A(n2174), .Z(n2008) );
  CIVX2 U1681 ( .A(reset), .Z(n2015) );
  CIVX2 U1682 ( .A(n2166), .Z(n2016) );
  CIVX2 U1697 ( .A(res_not_wire[62]), .Z(n2031) );
  CIVX2 U1708 ( .A(result[37]), .Z(n2042) );
  CIVX2 U1711 ( .A(result[41]), .Z(n2045) );
  CIVX2 U1717 ( .A(result[31]), .Z(n2051) );
  CIVX2 U1719 ( .A(result[29]), .Z(n2053) );
  CIVX2 U1734 ( .A(result[30]), .Z(n2068) );
  CIVX2 U1754 ( .A(res_not_wire[48]), .Z(n2088) );
  CIVX2 U1756 ( .A(res_not_wire[54]), .Z(n2090) );
  CIVX2 U1761 ( .A(res_not_wire[42]), .Z(n2095) );
  CIVX2 U1767 ( .A(n2255), .Z(n2101) );
  CIVX2 U1771 ( .A(n2227), .Z(n2105) );
  CIVX2 U1783 ( .A(n2222), .Z(n2117) );
  CIVX2 U1784 ( .A(n2217), .Z(n2118) );
  CIVX2 U1790 ( .A(res_not_wire[24]), .Z(n2124) );
  CIVX2 U1791 ( .A(res_not_wire[18]), .Z(n2125) );
  CIVX2 U1796 ( .A(n2212), .Z(n2130) );
  CIVX2 U1804 ( .A(res_not_wire[0]), .Z(n2138) );
  CIVX2 U1806 ( .A(n2834), .Z(n2140) );
  CIVX2 U1807 ( .A(n53), .Z(n2141) );
  CIVX2 U1809 ( .A(i[8]), .Z(n2143) );
  CIVX2 U1810 ( .A(n2207), .Z(n2144) );
  CIVX2 U1812 ( .A(n2195), .Z(n2146) );
  CIVX2 U1814 ( .A(n2190), .Z(n2148) );
  CIVX2 U1815 ( .A(n2185), .Z(n2149) );
  CIVX2 U1818 ( .A(n2180), .Z(n2150) );
  CIVX2 U1827 ( .A(n962), .Z(n2159) );
  CAOR2X1 U1832 ( .A(i[31]), .B(n2007), .C(n2169), .D(n3005), .Z(n955) );
  COR4X1 U1833 ( .A(n2155), .B(n2179), .C(i[5]), .D(n2180), .Z(n2175) );
  COR4X1 U1834 ( .A(n2163), .B(n2179), .C(i[7]), .D(n2185), .Z(n2189) );
  COR4X1 U1835 ( .A(n2143), .B(n2179), .C(i[9]), .D(n2190), .Z(n2194) );
  COR4X1 U1836 ( .A(n2154), .B(n2179), .C(i[11]), .D(n2195), .Z(n2199) );
  CND2IX1 U1837 ( .B(n2202), .A(i[12]), .Z(n2201) );
  COR4X1 U1838 ( .A(n2153), .B(n2179), .C(i[13]), .D(n2200), .Z(n2203) );
  COR4X1 U1839 ( .A(n2129), .B(n2179), .C(i[16]), .D(n2207), .Z(n2211) );
  COR4X1 U1840 ( .A(n2119), .B(n2179), .C(i[18]), .D(n2212), .Z(n2216) );
  COR4X1 U1841 ( .A(n2123), .B(n2179), .C(i[20]), .D(n2217), .Z(n2221) );
  COR4X1 U1842 ( .A(n2122), .B(n2179), .C(i[22]), .D(n2222), .Z(n2226) );
  CND2IX1 U1844 ( .B(n2234), .A(n2103), .Z(n2233) );
  COR4X1 U1845 ( .A(n2103), .B(n2179), .C(i[26]), .D(n2234), .Z(n2236) );
  COR4X1 U1846 ( .A(n2179), .B(n2102), .C(n2100), .D(i[28]), .Z(n2240) );
  CAOR2X1 U1847 ( .A(valid), .B(n2874), .C(n3004), .D(n3586), .Z(n923) );
  CAN4X1 U1848 ( .A(n2249), .B(n2252), .C(n2253), .D(n2254), .Z(n2166) );
  CAN4X1 U1874 ( .A(n56), .B(n53), .C(n1119), .D(reset), .Z(n2256) );
  CNR8X1 U1875 ( .A(i[1]), .B(i[19]), .C(i[16]), .D(i[2]), .E(n2839), .F(n2840), .G(n2837), .H(n2841), .Z(n2255) );
  COR3X1 U1876 ( .A(i[0]), .B(i[11]), .C(n2842), .Z(n2841) );
  COR6X1 U1877 ( .A(i[11]), .B(n2842), .C(n2840), .D(i[5]), .E(i[19]), .F(
        i[16]), .Z(n2843) );
  COR8X1 U1878 ( .A(i[20]), .B(i[17]), .C(i[22]), .D(i[21]), .E(i[26]), .F(
        i[24]), .G(i[9]), .H(i[30]), .Z(n2842) );
  COR8X1 U1879 ( .A(i[13]), .B(i[12]), .C(i[10]), .D(n2844), .E(i[28]), .F(
        i[27]), .G(i[25]), .H(n2845), .Z(n2840) );
  COR4X1 U1880 ( .A(i[29]), .B(i[6]), .C(i[7]), .D(i[8]), .Z(n2845) );
  COR4X1 U1881 ( .A(i[14]), .B(i[15]), .C(i[18]), .D(i[23]), .Z(n2844) );
  CND2IX1 U1882 ( .B(n2892), .A(nst[1]), .Z(n52) );
  CFD1XL \res_not_reg[54]  ( .D(n865), .CP(clock), .Q(res_not_wire[54]), .QN(
        n2960) );
  CFD1XL \res_not_reg[30]  ( .D(n889), .CP(clock), .Q(res_not_wire[30]), .QN(
        n2988) );
  CFD1QXL \result_reg[31]  ( .D(n794), .CP(clock), .Q(result[31]) );
  CFD1XL \res_not_reg[59]  ( .D(n860), .CP(clock), .Q(n2851), .QN(n106) );
  CFD1QXL \result_reg[29]  ( .D(n2891), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[30]  ( .D(n795), .CP(clock), .Q(result[30]) );
  CFD1XL \res_not_reg[55]  ( .D(n864), .CP(clock), .QN(n110) );
  CFD1XL \res_not_reg[51]  ( .D(n868), .CP(clock), .QN(n114) );
  CFD1XL \res_not_reg[53]  ( .D(n866), .CP(clock), .Q(n2888), .QN(n112) );
  CFD1XL \res_not_reg[49]  ( .D(n870), .CP(clock), .QN(n116) );
  CFD1XL \res_not_reg[33]  ( .D(n886), .CP(clock), .Q(n2965), .QN(n2852) );
  CFD1XL \res_not_reg[47]  ( .D(n872), .CP(clock), .QN(n118) );
  CFD1XL \res_not_reg[35]  ( .D(n884), .CP(clock), .QN(n130) );
  CFD1XL \res_not_reg[41]  ( .D(n878), .CP(clock), .Q(n2850), .QN(n124) );
  CFD1XL \res_not_reg[31]  ( .D(n888), .CP(clock), .Q(n2886), .QN(n134) );
  CFD1XL \res_not_reg[36]  ( .D(n883), .CP(clock), .Q(res_not_wire[36]), .QN(
        n2955) );
  CFD1XL \res_not_reg[37]  ( .D(n882), .CP(clock), .QN(n128) );
  CFD1XL \res_not_reg[43]  ( .D(n876), .CP(clock), .Q(n2848), .QN(n122) );
  CFD1XL \res_not_reg[23]  ( .D(n896), .CP(clock), .QN(n142) );
  CFD1XL \res_not_reg[25]  ( .D(n894), .CP(clock), .QN(n140) );
  CFD1XL \res_not_reg[29]  ( .D(n890), .CP(clock), .QN(n136) );
  CFD1XL \res_not_reg[27]  ( .D(n892), .CP(clock), .Q(n2856), .QN(n138) );
  CFD1XL \res_not_reg[45]  ( .D(n874), .CP(clock), .Q(n2887), .QN(n120) );
  CFD1XL \result_reg[49]  ( .D(n839), .CP(clock), .Q(result[49]), .QN(n2962)
         );
  CFD1XL \res_not_reg[21]  ( .D(n898), .CP(clock), .QN(n144) );
  CFD1XL \res_not_reg[17]  ( .D(n902), .CP(clock), .QN(n148) );
  CFD1XL \res_not_reg[19]  ( .D(n900), .CP(clock), .Q(n2885), .QN(n146) );
  CFD1XL \result_reg[48]  ( .D(n840), .CP(clock), .Q(result[48]), .QN(n2963)
         );
  CFD1XL \res_not_reg[11]  ( .D(n908), .CP(clock), .QN(n154) );
  CFD1XL \res_not_reg[15]  ( .D(n904), .CP(clock), .Q(n2884), .QN(n150) );
  CFD1XL \result_reg[38]  ( .D(n850), .CP(clock), .Q(result[38]), .QN(n2961)
         );
  CFD1XL \result_reg[39]  ( .D(n849), .CP(clock), .Q(result[39]), .QN(n2964)
         );
  CFD1XL \result_reg[40]  ( .D(n848), .CP(clock), .Q(result[40]), .QN(n2957)
         );
  CFD1XL \res_not_reg[4]  ( .D(n915), .CP(clock), .Q(res_not_wire[4]) );
  CFD1XL \res_not_reg[5]  ( .D(n914), .CP(clock), .QN(n160) );
  CFD1XL \res_not_reg[7]  ( .D(n912), .CP(clock), .Q(n2880), .QN(n158) );
  CTSX2 A2 ( .A(1'b0), .E(n2876), .Z(c_inop1) );
  CTSX2 A1 ( .A(1'b1), .E(opera1[31]), .Z(c_inop1) );
  CFD1XL \result_reg[35]  ( .D(n853), .CP(clock), .Q(result[35]), .QN(n2953)
         );
  CFD1XL \res_not_reg[3]  ( .D(n916), .CP(clock), .Q(n2854), .QN(n162) );
  CFD1XL \res_not_reg[0]  ( .D(n920), .CP(clock), .Q(res_not_wire[0]), .QN(
        n2937) );
  CFD1QXL \result_reg[63]  ( .D(n919), .CP(clock), .Q(result[63]) );
  CFD4QXL \cst_reg[0]  ( .D(n55), .CP(clock), .SD(n2015), .Q(n56) );
  CFD4QXL \cst_reg[1]  ( .D(n52), .CP(clock), .SD(n2015), .Q(n53) );
  CFD2XL \cst_reg[2]  ( .D(N34), .CP(clock), .CD(n2015), .Q(n3584), .QN(n1119)
         );
  CFD1XL \res_not_reg[39]  ( .D(n880), .CP(clock), .Q(n3165), .QN(n126) );
  CFD1X1 sign_reg ( .D(n2893), .CP(clock), .Q(n1061), .QN(n2137) );
  CFD1QXL valid_reg ( .D(n923), .CP(clock), .Q(valid) );
  CFD1QXL \i_reg[8]  ( .D(n946), .CP(clock), .Q(i[8]) );
  CFD1QXL \res_not_reg[38]  ( .D(n881), .CP(clock), .Q(res_not_wire[38]) );
  CFD1QXL \res_not_reg[32]  ( .D(n887), .CP(clock), .Q(res_not_wire[32]) );
  CFD1QXL \res_not_reg[2]  ( .D(n917), .CP(clock), .Q(res_not_wire[2]) );
  CFD1QXL \res_not_reg[14]  ( .D(n905), .CP(clock), .Q(res_not_wire[14]) );
  CFD1QXL \res_not_reg[13]  ( .D(n906), .CP(clock), .Q(n960) );
  CFD1QXL \res_not_reg[10]  ( .D(n909), .CP(clock), .Q(res_not_wire[10]) );
  CFD1QXL \res_not_reg[8]  ( .D(n911), .CP(clock), .Q(res_not_wire[8]) );
  CFD1QXL \res_not_reg[28]  ( .D(n891), .CP(clock), .Q(res_not_wire[28]) );
  CFD1QXL \res_not_reg[26]  ( .D(n893), .CP(clock), .Q(res_not_wire[26]) );
  CFD1QXL \res_not_reg[24]  ( .D(n895), .CP(clock), .Q(res_not_wire[24]) );
  CFD1QXL \res_not_reg[63]  ( .D(n793), .CP(clock), .Q(n1056) );
  CFD1QXL \res_not_reg[62]  ( .D(n857), .CP(clock), .Q(res_not_wire[62]) );
  CFD1QXL \res_not_reg[61]  ( .D(n858), .CP(clock), .Q(n1053) );
  CFD1QXL \res_not_reg[60]  ( .D(n859), .CP(clock), .Q(res_not_wire[60]) );
  CFD1QXL \res_not_reg[58]  ( .D(n861), .CP(clock), .Q(res_not_wire[58]) );
  CFD1QXL \res_not_reg[57]  ( .D(n862), .CP(clock), .Q(n1093) );
  CFD1QXL \res_not_reg[56]  ( .D(n863), .CP(clock), .Q(res_not_wire[56]) );
  CFD1QXL \res_not_reg[52]  ( .D(n867), .CP(clock), .Q(res_not_wire[52]) );
  CFD1QXL \res_not_reg[50]  ( .D(n869), .CP(clock), .Q(res_not_wire[50]) );
  CFD1QXL \res_not_reg[48]  ( .D(n871), .CP(clock), .Q(res_not_wire[48]) );
  CFD1QXL \res_not_reg[46]  ( .D(n873), .CP(clock), .Q(res_not_wire[46]) );
  CFD1QXL \res_not_reg[44]  ( .D(n875), .CP(clock), .Q(res_not_wire[44]) );
  CFD1QXL \res_not_reg[42]  ( .D(n877), .CP(clock), .Q(res_not_wire[42]) );
  CFD1QXL \res_not_reg[40]  ( .D(n879), .CP(clock), .Q(res_not_wire[40]) );
  CFD1QXL \res_not_reg[22]  ( .D(n897), .CP(clock), .Q(res_not_wire[22]) );
  CFD1QXL \res_not_reg[20]  ( .D(n899), .CP(clock), .Q(res_not_wire[20]) );
  CFD1QXL \res_not_reg[18]  ( .D(n901), .CP(clock), .Q(res_not_wire[18]) );
  CFD1QXL \res_not_reg[16]  ( .D(n903), .CP(clock), .Q(res_not_wire[16]) );
  CFD1QXL \res_not_reg[9]  ( .D(n910), .CP(clock), .Q(n962) );
  CFD1QXL \res_not_reg[6]  ( .D(n913), .CP(clock), .Q(res_not_wire[6]) );
  CFD1QXL \res_not_reg[34]  ( .D(n885), .CP(clock), .Q(res_not_wire[34]) );
  CFD1QXL \result_reg[47]  ( .D(n841), .CP(clock), .Q(result[47]) );
  CFD1QXL \result_reg[34]  ( .D(n854), .CP(clock), .Q(result[34]) );
  CFD1QXL \result_reg[36]  ( .D(n852), .CP(clock), .Q(result[36]) );
  CFD1QXL \result_reg[41]  ( .D(n847), .CP(clock), .Q(result[41]) );
  CFD1QXL \result_reg[52]  ( .D(n836), .CP(clock), .Q(result[52]) );
  CFD1QXL \result_reg[46]  ( .D(n842), .CP(clock), .Q(result[46]) );
  CFD1QXL \result_reg[37]  ( .D(n851), .CP(clock), .Q(result[37]) );
  CFD1QXL \result_reg[50]  ( .D(n838), .CP(clock), .Q(result[50]) );
  CFD1QXL \result_reg[42]  ( .D(n846), .CP(clock), .Q(result[42]) );
  CFD1QXL \result_reg[43]  ( .D(n845), .CP(clock), .Q(result[43]) );
  CFD1QXL \result_reg[51]  ( .D(n837), .CP(clock), .Q(result[51]) );
  CFD1QXL \result_reg[53]  ( .D(n835), .CP(clock), .Q(result[53]) );
  CFD1QXL \result_reg[54]  ( .D(n834), .CP(clock), .Q(result[54]) );
  CFD1QXL \result_reg[44]  ( .D(n844), .CP(clock), .Q(result[44]) );
  CFD1QXL \result_reg[57]  ( .D(n831), .CP(clock), .Q(result[57]) );
  CFD1QXL \result_reg[45]  ( .D(n843), .CP(clock), .Q(result[45]) );
  CFD1QXL \result_reg[55]  ( .D(n833), .CP(clock), .Q(result[55]) );
  CFD1QXL \result_reg[56]  ( .D(n832), .CP(clock), .Q(result[56]) );
  CFD1QXL \result_reg[59]  ( .D(n829), .CP(clock), .Q(result[59]) );
  CFD1QXL \result_reg[58]  ( .D(n830), .CP(clock), .Q(result[58]) );
  CFD1QXL \result_reg[60]  ( .D(n828), .CP(clock), .Q(result[60]) );
  CFD1XL \nst_reg[1]  ( .D(n2894), .CP(clock), .Q(nst[1]), .QN(n2049) );
  CFD1XL \nst_reg[2]  ( .D(n921), .CP(clock), .Q(nst[2]) );
  CFD1XL \nst_reg[0]  ( .D(n2896), .CP(clock), .Q(nst[0]) );
  CFD1XL \i_reg[0]  ( .D(n952), .CP(clock), .Q(i[0]), .QN(n2162) );
  CFD1XL \i_reg[1]  ( .D(n951), .CP(clock), .Q(i[1]), .QN(n2157) );
  CFD1XL \i_reg[23]  ( .D(n931), .CP(clock), .Q(i[23]), .QN(n2106) );
  CFD1XL \i_reg[21]  ( .D(n933), .CP(clock), .Q(i[21]), .QN(n2122) );
  CFD1XL \i_reg[19]  ( .D(n935), .CP(clock), .Q(i[19]), .QN(n2123) );
  CFD1XL \i_reg[17]  ( .D(n937), .CP(clock), .Q(i[17]), .QN(n2119) );
  CFD1XL \i_reg[15]  ( .D(n939), .CP(clock), .Q(i[15]), .QN(n2129) );
  CFD1XL \i_reg[10]  ( .D(n944), .CP(clock), .Q(i[10]), .QN(n2154) );
  CFD1XL \i_reg[4]  ( .D(n949), .CP(clock), .Q(i[4]), .QN(n2155) );
  CFD1XL \i_reg[25]  ( .D(n929), .CP(clock), .Q(i[25]), .QN(n2103) );
  CFD1XL \i_reg[22]  ( .D(n932), .CP(clock), .Q(i[22]) );
  CFD1XL \i_reg[7]  ( .D(n947), .CP(clock), .Q(i[7]) );
  CFD1XL \i_reg[6]  ( .D(n948), .CP(clock), .Q(i[6]), .QN(n2163) );
  CFD1XL \i_reg[27]  ( .D(n927), .CP(clock), .Q(i[27]), .QN(n2102) );
  CFD1XL \i_reg[20]  ( .D(n934), .CP(clock), .Q(i[20]) );
  CFD1XL \i_reg[18]  ( .D(n936), .CP(clock), .Q(i[18]) );
  CFD1XL \i_reg[9]  ( .D(n945), .CP(clock), .Q(i[9]) );
  CFD1XL \i_reg[5]  ( .D(n953), .CP(clock), .Q(i[5]) );
  CFD1XL \i_reg[16]  ( .D(n938), .CP(clock), .Q(i[16]) );
  CFD1XL \i_reg[11]  ( .D(n943), .CP(clock), .Q(i[11]) );
  CFD1XL \i_reg[26]  ( .D(n928), .CP(clock), .Q(i[26]), .QN(n2121) );
  CFD1XL \i_reg[3]  ( .D(n954), .CP(clock), .Q(i[3]), .QN(n2151) );
  CFD1XL \i_reg[24]  ( .D(n930), .CP(clock), .Q(i[24]), .QN(n2863) );
  CFD1XL \i_reg[28]  ( .D(n926), .CP(clock), .Q(i[28]) );
  CFD1XL \i_reg[31]  ( .D(n955), .CP(clock), .Q(i[31]), .QN(n2847) );
  CFD1XL \i_reg[12]  ( .D(n942), .CP(clock), .Q(i[12]), .QN(n2153) );
  CFD1XL \i_reg[2]  ( .D(n950), .CP(clock), .Q(i[2]), .QN(n2156) );
  CFD1XL \i_reg[29]  ( .D(n925), .CP(clock), .Q(i[29]), .QN(n2120) );
  CFD1XL \i_reg[30]  ( .D(n2898), .CP(clock), .Q(i[30]), .QN(n2104) );
  CFD1XL \i_reg[13]  ( .D(n941), .CP(clock), .Q(i[13]), .QN(n2152) );
  CFD1XL \i_reg[14]  ( .D(n940), .CP(clock), .Q(i[14]) );
  CFD1XL \res_not_reg[12]  ( .D(n907), .CP(clock), .Q(res_not_wire[12]), .QN(
        n2147) );
  CFD1XL \result_reg[23]  ( .D(n802), .CP(clock), .Q(result[23]), .QN(n2056)
         );
  CFD1XL \result_reg[26]  ( .D(n2899), .CP(clock), .Q(result[26]), .QN(n2070)
         );
  CFD1XL \result_reg[14]  ( .D(n811), .CP(clock), .Q(result[14]), .QN(n2076)
         );
  CFD1XL \result_reg[27]  ( .D(n798), .CP(clock), .Q(result[27]), .QN(n2054)
         );
  CFD1XL \result_reg[20]  ( .D(n805), .CP(clock), .Q(result[20]), .QN(n2073)
         );
  CFD1XL \result_reg[17]  ( .D(n808), .CP(clock), .Q(result[17]), .QN(n2059)
         );
  CFD1XL \result_reg[11]  ( .D(n814), .CP(clock), .Q(result[11]), .QN(n2062)
         );
  CFD1XL \result_reg[8]  ( .D(n817), .CP(clock), .Q(result[8]), .QN(n2079) );
  CFD1XL \result_reg[5]  ( .D(n820), .CP(clock), .Q(result[5]), .QN(n2065) );
  CFD1XL \result_reg[2]  ( .D(n823), .CP(clock), .Q(result[2]), .QN(n2081) );
  CFD1XL \result_reg[25]  ( .D(n2900), .CP(clock), .Q(result[25]), .QN(n2055)
         );
  CFD1XL \result_reg[22]  ( .D(n803), .CP(clock), .Q(result[22]), .QN(n2072)
         );
  CFD1XL \result_reg[18]  ( .D(n807), .CP(clock), .Q(result[18]), .QN(n2074)
         );
  CFD1XL \result_reg[16]  ( .D(n809), .CP(clock), .Q(result[16]), .QN(n2075)
         );
  CFD1XL \result_reg[15]  ( .D(n810), .CP(clock), .Q(result[15]), .QN(n2060)
         );
  CFD1XL \result_reg[13]  ( .D(n812), .CP(clock), .Q(result[13]), .QN(n2061)
         );
  CFD1XL \result_reg[12]  ( .D(n2904), .CP(clock), .Q(result[12]), .QN(n2077)
         );
  CFD1XL \result_reg[10]  ( .D(n815), .CP(clock), .Q(result[10]), .QN(n2078)
         );
  CFD1XL \result_reg[9]  ( .D(n2906), .CP(clock), .Q(result[9]), .QN(n2063) );
  CFD1XL \result_reg[7]  ( .D(n818), .CP(clock), .Q(result[7]), .QN(n2064) );
  CFD1XL \result_reg[6]  ( .D(n819), .CP(clock), .Q(result[6]), .QN(n2052) );
  CFD1XL \result_reg[4]  ( .D(n821), .CP(clock), .Q(result[4]), .QN(n2080) );
  CFD1XL \result_reg[3]  ( .D(n822), .CP(clock), .Q(result[3]), .QN(n2066) );
  CFD1XL \result_reg[1]  ( .D(n824), .CP(clock), .Q(result[1]), .QN(n2067) );
  CFD1XL \result_reg[0]  ( .D(n2908), .CP(clock), .Q(result[0]), .QN(n3579) );
  CFD1XL \result_reg[19]  ( .D(n2909), .CP(clock), .Q(result[19]), .QN(n2058)
         );
  CFD1XL \result_reg[24]  ( .D(n2910), .CP(clock), .Q(result[24]), .QN(n2071)
         );
  CFD1XL \result_reg[21]  ( .D(n2911), .CP(clock), .Q(result[21]), .QN(n2057)
         );
  CFD1XL \result_reg[28]  ( .D(n797), .CP(clock), .Q(result[28]), .QN(n2069)
         );
  CFD1XL \res_not_reg[1]  ( .D(n918), .CP(clock), .QN(n164) );
  CFD1QXL \result_reg[62]  ( .D(n826), .CP(clock), .Q(result[62]) );
  CFD1XL \result_reg[32]  ( .D(n2912), .CP(clock), .Q(result[32]) );
  CFD1XL \result_reg[33]  ( .D(n855), .CP(clock), .Q(result[33]), .QN(n2928)
         );
  CFD1QXL \result_reg[61]  ( .D(n827), .CP(clock), .Q(result[61]) );
  COND11X1 U1883 ( .A(n2179), .B(i[1]), .C(n2162), .D(n2181), .Z(n951) );
  CNR2IX1 U1884 ( .B(result[32]), .A(n3001), .Z(n3159) );
  CND2X2 U1885 ( .A(n3198), .B(n3197), .Z(n3205) );
  CANR4CX2 U1886 ( .A(n3180), .B(n3417), .C(n3181), .D(n3456), .Z(n3186) );
  CENX2 U1887 ( .A(result[36]), .B(n2846), .Z(n3180) );
  CNIVX1 U1888 ( .A(n3135), .Z(n2846) );
  COND1X1 U1889 ( .A(n3167), .B(n3166), .C(n3173), .Z(n3171) );
  CND2X2 U1890 ( .A(n3167), .B(n3166), .Z(n3173) );
  CND2XL U1891 ( .A(n3355), .B(res_not_wire[58]), .Z(n3560) );
  CND2X2 U1892 ( .A(result[0]), .B(n3574), .Z(n3558) );
  CANR1X1 U1893 ( .A(n3437), .B(n3208), .C(n3207), .Z(n3447) );
  CANR1X1 U1894 ( .A(n3242), .B(n3255), .C(n3241), .Z(n3486) );
  CND2IXL U1895 ( .B(n3018), .A(n2927), .Z(n3161) );
  CENX1 U1896 ( .A(n2138), .B(c_inres), .Z(n2634) );
  CENX1 U1897 ( .A(n3512), .B(n3511), .Z(n3513) );
  CND2IX1 U1898 ( .B(n3501), .A(n2932), .Z(n3314) );
  CENX1 U1899 ( .A(res_not_wire[28]), .B(n3021), .Z(n3022) );
  CENX1 U1900 ( .A(n106), .B(n3560), .Z(n3402) );
  CEOX1 U1901 ( .A(opera1[6]), .B(opera1[31]), .Z(n3166) );
  COR2X1 U1902 ( .A(n3380), .B(n3364), .Z(n3386) );
  CND2X1 U1903 ( .A(n2847), .B(n2843), .Z(n2837) );
  CND3XL U1904 ( .A(n3058), .B(res_not_wire[16]), .C(n2884), .Z(n3050) );
  CNR2X1 U1905 ( .A(n2116), .B(n130), .Z(n3130) );
  CNR2IX1 U1906 ( .B(res_not_wire[52]), .A(n3314), .Z(n2997) );
  COND3X1 U1907 ( .A(n2852), .B(n3161), .C(n2869), .D(n3122), .Z(n3129) );
  CND2IX1 U1908 ( .B(n3235), .A(n3227), .Z(n3236) );
  CEOX1 U1909 ( .A(opera1[16]), .B(opera1[31]), .Z(n3229) );
  CEOX1 U1910 ( .A(opera1[8]), .B(opera1[31]), .Z(n3168) );
  COR2X1 U1911 ( .A(n148), .B(n3050), .Z(n3052) );
  CENX1 U1912 ( .A(n3368), .B(n3367), .Z(n3373) );
  CND2X1 U1913 ( .A(res_not_wire[46]), .B(n2994), .Z(n3262) );
  CMXI2XL U1914 ( .A0(n3410), .A1(n3409), .S(result[32]), .Z(n3411) );
  CND3XL U1915 ( .A(n2644), .B(n3101), .C(n3100), .Z(n823) );
  CNR2XL U1916 ( .A(n2034), .B(n3553), .Z(n3533) );
  COND1XL U1917 ( .A(n3230), .B(n3229), .C(n3246), .Z(n3243) );
  CENX1 U1918 ( .A(n3380), .B(n3364), .Z(n3384) );
  COAN1X1 U1919 ( .A(n3177), .B(n3176), .C(n3204), .Z(n3179) );
  CND2IX1 U1920 ( .B(n3143), .A(result[37]), .Z(n3454) );
  CND2X1 U1921 ( .A(n2854), .B(n3094), .Z(n3092) );
  CND2X1 U1922 ( .A(n3013), .B(n962), .Z(n3014) );
  CND2X1 U1923 ( .A(n2986), .B(n2875), .Z(n3044) );
  CND2XL U1924 ( .A(n2834), .B(n3553), .Z(n3035) );
  CND2X1 U1925 ( .A(n2852), .B(n3161), .Z(n3122) );
  CND2X1 U1926 ( .A(n2955), .B(n3416), .Z(n3146) );
  CEOX1 U1927 ( .A(n3540), .B(n3539), .Z(n2853) );
  CEOX1 U1928 ( .A(opera1[9]), .B(opera1[31]), .Z(n3176) );
  CND2X1 U1929 ( .A(n3211), .B(n3210), .Z(n3218) );
  CIVX1 U1930 ( .A(n3212), .Z(n3211) );
  CNR2X1 U1931 ( .A(n3173), .B(n3172), .Z(n3169) );
  CENX1 U1932 ( .A(n3290), .B(n3289), .Z(n3291) );
  COR2X1 U1933 ( .A(n3086), .B(n160), .Z(n3088) );
  CND3XL U1934 ( .A(n3013), .B(n962), .C(res_not_wire[10]), .Z(n3068) );
  CNR2IX1 U1935 ( .B(res_not_wire[18]), .A(n3052), .Z(n2986) );
  CND8X1 U1936 ( .A(n2848), .B(n2849), .C(n2850), .D(n2887), .E(
        res_not_wire[36]), .F(res_not_wire[44]), .G(res_not_wire[42]), .H(
        res_not_wire[40]), .Z(n2995) );
  CIVX2 U1937 ( .A(n3225), .Z(n2849) );
  CND2X1 U1938 ( .A(n3454), .B(n3144), .Z(n3456) );
  COND1XL U1939 ( .A(n3142), .B(n3105), .C(n3115), .Z(n3112) );
  CIVX1 U1940 ( .A(n3109), .Z(n3142) );
  CND2X1 U1941 ( .A(i[30]), .B(i[29]), .Z(n3007) );
  CND4X1 U1942 ( .A(n2851), .B(n3355), .C(res_not_wire[58]), .D(
        res_not_wire[60]), .Z(n3562) );
  CNR2X1 U1943 ( .A(n2852), .B(n3161), .Z(n2933) );
  COND3XL U1944 ( .A(n2853), .B(n3558), .C(n3543), .D(n3542), .Z(n831) );
  CEOX1 U1945 ( .A(opera1[13]), .B(opera1[31]), .Z(n3216) );
  COND1XL U1946 ( .A(n3200), .B(n3199), .C(n3212), .Z(n3209) );
  COND1XL U1947 ( .A(n3169), .B(n3168), .C(n3178), .Z(n3175) );
  CND3X1 U1948 ( .A(res_not_wire[4]), .B(n2854), .C(n3094), .Z(n3086) );
  CND2XL U1949 ( .A(n3031), .B(res_not_wire[24]), .Z(n3029) );
  CIVX2 U1950 ( .A(n3033), .Z(n3031) );
  CNR2X1 U1951 ( .A(n2960), .B(n110), .Z(n2991) );
  COND2X1 U1952 ( .A(n3299), .B(n2097), .C(n3495), .D(n3494), .Z(n2855) );
  CIVX1 U1953 ( .A(n2855), .Z(n3308) );
  CND2X1 U1954 ( .A(n2928), .B(n3154), .Z(n3110) );
  CENX1 U1955 ( .A(n3115), .B(n3138), .Z(n3131) );
  CND2X1 U1956 ( .A(n2856), .B(n3023), .Z(n3021) );
  CIVXL U1957 ( .A(n3025), .Z(n3023) );
  CNR2X1 U1958 ( .A(n144), .B(n3044), .Z(n2952) );
  CAN4X1 U1959 ( .A(n2939), .B(n2965), .C(n2927), .D(n2857), .Z(n2994) );
  CIVX1 U1960 ( .A(n3018), .Z(n2857) );
  CNR3XL U1961 ( .A(n3581), .B(n114), .C(n116), .Z(n2932) );
  CND3XL U1962 ( .A(n2682), .B(n3082), .C(n3081), .Z(n817) );
  CEOXL U1963 ( .A(n2954), .B(n128), .Z(n3472) );
  CEOXL U1964 ( .A(n1053), .B(n3562), .Z(n3552) );
  CEOX1 U1965 ( .A(opera1[12]), .B(opera1[31]), .Z(n3210) );
  CEOX1 U1966 ( .A(opera1[10]), .B(opera1[31]), .Z(n3197) );
  CND2IX1 U1967 ( .B(n3246), .A(n3244), .Z(n3290) );
  CND2X1 U1968 ( .A(n3233), .B(n3232), .Z(n2864) );
  CENX1 U1969 ( .A(n3173), .B(n3172), .Z(n3174) );
  CEOX1 U1970 ( .A(opera1[0]), .B(opera1[31]), .Z(n2958) );
  CND2IX1 U1971 ( .B(n3088), .A(res_not_wire[6]), .Z(n3077) );
  COR2X1 U1972 ( .A(n154), .B(n3068), .Z(n3070) );
  COR2X1 U1973 ( .A(n142), .B(n3034), .Z(n3033) );
  COND1XL U1974 ( .A(n3339), .B(n3338), .C(n3368), .Z(n3372) );
  COND2X1 U1975 ( .A(n2953), .B(n3131), .C(n3133), .D(n3132), .Z(n2858) );
  CIVX2 U1976 ( .A(n2858), .Z(n3417) );
  CENX1 U1977 ( .A(res_not_wire[4]), .B(n3092), .Z(n3093) );
  CND2X1 U1978 ( .A(n3058), .B(n2884), .Z(n3056) );
  CENX1 U1979 ( .A(n3052), .B(res_not_wire[18]), .Z(n3049) );
  CND2X1 U1980 ( .A(n2989), .B(n2991), .Z(n2984) );
  COR2X1 U1981 ( .A(n118), .B(n3262), .Z(n3226) );
  COR4X1 U1982 ( .A(n138), .B(n136), .C(n2859), .D(n3025), .Z(n3018) );
  CIVX2 U1983 ( .A(res_not_wire[28]), .Z(n2859) );
  CND3XL U1984 ( .A(n2758), .B(n3047), .C(n3046), .Z(n805) );
  CND2IXL U1985 ( .B(n3558), .A(n3547), .Z(n3550) );
  COR3X1 U1986 ( .A(n3317), .B(n3323), .C(n3322), .Z(n3333) );
  COND1XL U1987 ( .A(n3211), .B(n3210), .C(n3218), .Z(n3213) );
  CENX1 U1988 ( .A(n3235), .B(n3234), .Z(n3240) );
  COND1XL U1989 ( .A(n3198), .B(n3197), .C(n3205), .Z(n3206) );
  CND2IX1 U1990 ( .B(opera2[0]), .A(opera2_63), .Z(n2948) );
  CND4X1 U1991 ( .A(n3028), .B(res_not_wire[26]), .C(res_not_wire[24]), .D(
        n3031), .Z(n3025) );
  CANR1XL U1992 ( .A(n3504), .B(n3503), .C(n3502), .Z(n3293) );
  CEOX1 U1993 ( .A(result[62]), .B(n3385), .Z(n2946) );
  CND2XL U1994 ( .A(n160), .B(n3086), .Z(n3087) );
  CND2XL U1995 ( .A(n154), .B(n3068), .Z(n3069) );
  CND2XL U1996 ( .A(n148), .B(n3050), .Z(n3051) );
  CND4X1 U1997 ( .A(n3040), .B(n2986), .C(n2875), .D(res_not_wire[22]), .Z(
        n3034) );
  CNR3X1 U1998 ( .A(n2153), .B(n2200), .C(n2152), .Z(n2206) );
  CND3X1 U1999 ( .A(n2105), .B(i[23]), .C(i[24]), .Z(n2234) );
  CND2X1 U2000 ( .A(n2869), .B(n3473), .Z(n3463) );
  CND2XL U2001 ( .A(n2988), .B(n3018), .Z(n3016) );
  CND2IX1 U2002 ( .B(n3236), .A(n3228), .Z(n3233) );
  CENX1 U2003 ( .A(n3325), .B(n3317), .Z(n3329) );
  COND1XL U2004 ( .A(n3217), .B(n3216), .C(n3235), .Z(n3239) );
  COND1XL U2005 ( .A(n3179), .B(result[41]), .C(n3202), .Z(n3188) );
  CEOXL U2006 ( .A(n3044), .B(n144), .Z(n3041) );
  CND3X1 U2007 ( .A(n2146), .B(i[10]), .C(i[11]), .Z(n2200) );
  CND4X1 U2008 ( .A(n2989), .B(n2991), .C(n1093), .D(res_not_wire[56]), .Z(
        n3538) );
  CND2XL U2009 ( .A(n2960), .B(n3518), .Z(n3519) );
  CND2XL U2010 ( .A(n118), .B(n3262), .Z(n3263) );
  COAN1X1 U2011 ( .A(n3466), .B(n2860), .C(n3457), .Z(n3458) );
  CIVX2 U2012 ( .A(n3467), .Z(n2860) );
  COAN1X1 U2013 ( .A(n3503), .B(n2861), .C(n3504), .Z(n2940) );
  CIVX2 U2014 ( .A(n3505), .Z(n2861) );
  COND1XL U2015 ( .A(n2862), .B(n3021), .C(n136), .Z(n3019) );
  CIVX2 U2016 ( .A(res_not_wire[28]), .Z(n2862) );
  CND3XL U2017 ( .A(n2663), .B(n3091), .C(n3090), .Z(n820) );
  CND3XL U2018 ( .A(n2701), .B(n3073), .C(n3072), .Z(n814) );
  CND3XL U2019 ( .A(n2739), .B(n3055), .C(n3054), .Z(n808) );
  CND2XL U2020 ( .A(n142), .B(n3034), .Z(n3037) );
  CND2X1 U2021 ( .A(n2863), .B(n2105), .Z(n2230) );
  CEOXL U2022 ( .A(n3314), .B(res_not_wire[52]), .Z(n3305) );
  CEOX1 U2023 ( .A(n3132), .B(n3133), .Z(n3116) );
  CMXI2X2 U2024 ( .A0(n2137), .A1(n3121), .S(n2167), .Z(n2893) );
  COND1XL U2025 ( .A(n2051), .B(n3553), .C(n3411), .Z(n3414) );
  CND2IX1 U2026 ( .B(n3011), .A(n3010), .Z(n3553) );
  COND3X1 U2027 ( .A(n3395), .B(n3394), .C(n3393), .D(n3392), .Z(n826) );
  CND2IX1 U2028 ( .B(n2998), .A(n3403), .Z(n3394) );
  CANR1X2 U2029 ( .A(n3512), .B(n3328), .C(n3327), .Z(n3522) );
  COND2X2 U2030 ( .A(n3321), .B(n2036), .C(n3320), .D(n3319), .Z(n3512) );
  CENXL U2031 ( .A(n3397), .B(n3396), .Z(n3398) );
  CANR1X2 U2032 ( .A(n3397), .B(n3383), .C(n3382), .Z(n3555) );
  COND2X2 U2033 ( .A(n3376), .B(n2086), .C(n3529), .D(n3528), .Z(n3397) );
  CANR3X2 U2034 ( .A(n3389), .B(n3546), .C(n3388), .D(n3387), .Z(n3390) );
  CEOXL U2035 ( .A(n3505), .B(n3503), .Z(n2950) );
  COND2X2 U2036 ( .A(n3209), .B(n2046), .C(n3447), .D(n3446), .Z(n3427) );
  COND2X2 U2037 ( .A(n3300), .B(n2098), .C(n3308), .D(n3307), .Z(n3318) );
  COND2X2 U2038 ( .A(n2864), .B(n2112), .C(n3486), .D(n3485), .Z(n3266) );
  CND2X1 U2039 ( .A(n3169), .B(n3168), .Z(n3178) );
  CND3X1 U2040 ( .A(c_inop1), .B(n2930), .C(n2958), .Z(n3109) );
  CEOX1 U2041 ( .A(opera1[31]), .B(opera1[1]), .Z(n2930) );
  CND2X1 U2042 ( .A(result[32]), .B(n3406), .Z(n3153) );
  CND2X1 U2043 ( .A(c_inop2), .B(n2635), .Z(n2643) );
  CIVX2 U2044 ( .A(n3077), .Z(n3083) );
  CIVX2 U2045 ( .A(n3070), .Z(n3066) );
  CANR1X1 U2046 ( .A(n3349), .B(n3337), .C(n3336), .Z(n3370) );
  CNIVX1 U2047 ( .A(n3553), .Z(n3001) );
  CNIVX1 U2048 ( .A(n3553), .Z(n3000) );
  COND1XL U2049 ( .A(n2958), .B(c_inop1), .C(n3107), .Z(n3407) );
  CIVX2 U2050 ( .A(n3063), .Z(n3058) );
  COND1X1 U2051 ( .A(n3007), .B(n2246), .C(i[31]), .Z(n3009) );
  CND2X1 U2052 ( .A(i[14]), .B(n2206), .Z(n2207) );
  CENX1 U2053 ( .A(n3320), .B(n3318), .Z(n3301) );
  CENX1 U2054 ( .A(n3266), .B(n3265), .Z(n3267) );
  CENX1 U2055 ( .A(n2992), .B(n3347), .Z(n3354) );
  CIVX1 U2056 ( .A(n3553), .Z(n2871) );
  CIVDX1 U2057 ( .A(n3551), .Z0(n2867), .Z1(n2868) );
  CIVX3 U2058 ( .A(opera2_63), .Z(n2866) );
  CANR1X1 U2059 ( .A(n3427), .B(n3215), .C(n3214), .Z(n3237) );
  CND2IX2 U2060 ( .B(n2996), .A(n2981), .Z(n3063) );
  CND2X1 U2061 ( .A(c_inop1), .B(n2958), .Z(n3107) );
  CND3X2 U2062 ( .A(n2980), .B(res_not_wire[2]), .C(n3102), .Z(n3098) );
  CAN3XL U2063 ( .A(result[33]), .B(n3109), .C(n3108), .Z(n2879) );
  CND2X2 U2064 ( .A(n3083), .B(n2873), .Z(n3079) );
  CNR3X2 U2065 ( .A(n2103), .B(n2234), .C(n2121), .Z(n2241) );
  CND3X1 U2066 ( .A(i[27]), .B(n2241), .C(i[28]), .Z(n2246) );
  CIVDX1 U2067 ( .A(n2999), .Z0(n2869), .Z1(n2870) );
  CND2IXL U2068 ( .B(n3015), .A(n3553), .Z(n2998) );
  CND2IXL U2069 ( .B(n3015), .A(n3553), .Z(n3551) );
  CND2IX1 U2070 ( .B(n3015), .A(n3553), .Z(n2999) );
  CIVXL U2071 ( .A(n2206), .Z(n2145) );
  CND2X1 U2072 ( .A(n3359), .B(n3358), .Z(n3369) );
  CND2X1 U2073 ( .A(n3275), .B(n3274), .Z(n3296) );
  CND2X1 U2074 ( .A(n3339), .B(n3338), .Z(n3368) );
  CND2X1 U2075 ( .A(n3280), .B(n3279), .Z(n3323) );
  CND2X1 U2076 ( .A(n3361), .B(n3360), .Z(n3378) );
  CND2X1 U2077 ( .A(n3230), .B(n3229), .Z(n3246) );
  CND2IX1 U2078 ( .B(n3265), .A(n3266), .Z(n3287) );
  CEOX1 U2079 ( .A(result[61]), .B(n3384), .Z(n3556) );
  CEOX1 U2080 ( .A(result[60]), .B(n3381), .Z(n3396) );
  CEOX1 U2081 ( .A(result[57]), .B(n3372), .Z(n3371) );
  CEOX1 U2082 ( .A(result[58]), .B(n3373), .Z(n3539) );
  CEOX1 U2083 ( .A(result[55]), .B(n3329), .Z(n3521) );
  CEOX1 U2084 ( .A(result[52]), .B(n3300), .Z(n3307) );
  CEOX1 U2085 ( .A(result[47]), .B(n2864), .Z(n3485) );
  CEOX1 U2086 ( .A(result[53]), .B(n3321), .Z(n3320) );
  CEOX1 U2087 ( .A(result[38]), .B(n3171), .Z(n3466) );
  CEOX1 U2088 ( .A(result[50]), .B(n3291), .Z(n3502) );
  CND2X1 U2089 ( .A(n3316), .B(n3315), .Z(n3325) );
  CND2X1 U2090 ( .A(n3200), .B(n3199), .Z(n3212) );
  CND2X1 U2091 ( .A(n3278), .B(n3277), .Z(n3285) );
  CND2X1 U2092 ( .A(n3177), .B(n3176), .Z(n3204) );
  CND3XL U2093 ( .A(n3142), .B(n3141), .C(n3140), .Z(n3170) );
  CND2X1 U2094 ( .A(n3217), .B(n3216), .Z(n3235) );
  CND2X1 U2095 ( .A(n3331), .B(n3330), .Z(n3341) );
  CND2X1 U2096 ( .A(n3298), .B(n3297), .Z(n3299) );
  CND2X1 U2097 ( .A(n3363), .B(n3362), .Z(n3380) );
  CNIVXL U2098 ( .A(n2643), .Z(n2926) );
  CENX1 U2099 ( .A(opera2[2]), .B(opera2_63), .Z(n2649) );
  CENX1 U2100 ( .A(opera2[25]), .B(opera2_63), .Z(n2795) );
  CANR1X1 U2101 ( .A(n3375), .B(n2934), .C(n3374), .Z(n3529) );
  CEOX1 U2102 ( .A(result[59]), .B(n3376), .Z(n3528) );
  CANR2X1 U2103 ( .A(n3294), .B(n3293), .C(result[50]), .D(n3292), .Z(n3495)
         );
  CND3XL U2104 ( .A(n3288), .B(n3504), .C(n3287), .Z(n3294) );
  CEOX1 U2105 ( .A(result[51]), .B(n3299), .Z(n3494) );
  CEOX1 U2106 ( .A(result[48]), .B(n3243), .Z(n3265) );
  COND1X1 U2107 ( .A(n2879), .B(n3111), .C(n3110), .Z(n3123) );
  CNR3XL U2108 ( .A(n2157), .B(n2162), .C(n2156), .Z(n2173) );
  CND3XL U2109 ( .A(i[4]), .B(n2150), .C(i[5]), .Z(n2185) );
  CND2X1 U2110 ( .A(i[3]), .B(n2173), .Z(n2180) );
  CND3XL U2111 ( .A(i[8]), .B(n2148), .C(i[9]), .Z(n2195) );
  CND3XL U2112 ( .A(i[15]), .B(n2144), .C(i[16]), .Z(n2212) );
  CND3XL U2113 ( .A(i[17]), .B(n2130), .C(i[18]), .Z(n2217) );
  CND3XL U2114 ( .A(i[19]), .B(n2118), .C(i[20]), .Z(n2222) );
  CND3XL U2115 ( .A(i[21]), .B(n2117), .C(i[22]), .Z(n2227) );
  CENX1 U2116 ( .A(n3349), .B(n3348), .Z(n3350) );
  CEOX1 U2117 ( .A(result[35]), .B(n3131), .Z(n3133) );
  CND3XL U2118 ( .A(i[6]), .B(n2149), .C(i[7]), .Z(n2190) );
  CANR1XL U2119 ( .A(n3187), .B(n3189), .C(n3188), .Z(n3185) );
  CND3XL U2120 ( .A(n3187), .B(n3183), .C(n2951), .Z(n3184) );
  CANR1XL U2121 ( .A(n3038), .B(n3037), .C(n3036), .Z(n2778) );
  CNIVX2 U2122 ( .A(n957), .Z(n2896) );
  CENX1 U2123 ( .A(n2984), .B(n3587), .Z(n3346) );
  CND3XL U2124 ( .A(n3527), .B(n3526), .C(n3525), .Z(n834) );
  CENX1 U2125 ( .A(n2979), .B(n3306), .Z(n3313) );
  CND3XL U2126 ( .A(n3452), .B(n3451), .C(n3450), .Z(n846) );
  CENX1 U2127 ( .A(res_not_wire[46]), .B(n2994), .Z(n3491) );
  CENX1 U2128 ( .A(n116), .B(n3501), .Z(n3510) );
  CND2X1 U2129 ( .A(n2802), .B(n2807), .Z(n2813) );
  CAN2X1 U2130 ( .A(res_not_wire[8]), .B(n2880), .Z(n2873) );
  COAN1X1 U2131 ( .A(n2250), .B(n2101), .C(n3008), .Z(n2874) );
  CAN2X1 U2132 ( .A(res_not_wire[20]), .B(n2885), .Z(n2875) );
  CIVDX1 U2133 ( .A(opera1[31]), .Z0(n2876), .Z1(n2877) );
  COR2X1 U2134 ( .A(n2662), .B(n2668), .Z(n2878) );
  CAN2X1 U2135 ( .A(n2722), .B(n3573), .Z(n2881) );
  CEOX1 U2136 ( .A(opera1[5]), .B(opera1[31]), .Z(n2882) );
  COR2X1 U2137 ( .A(n2744), .B(n2738), .Z(n2883) );
  CND2X1 U2138 ( .A(n2947), .B(n2948), .Z(n2635) );
  CIVXL U2139 ( .A(opera2[30]), .Z(n2003) );
  CIVDX1 U2140 ( .A(n2942), .Z1(n2890) );
  CIVXL U2141 ( .A(opera2[31]), .Z(n2942) );
  CENXL U2142 ( .A(n2890), .B(n2833), .Z(n2829) );
  CND2IXL U2143 ( .B(n3414), .A(n3413), .Z(n794) );
  CNIVX1 U2144 ( .A(n796), .Z(n2891) );
  CEOXL U2145 ( .A(opera2[29]), .B(n2866), .Z(n2820) );
  CDLY1XL U2146 ( .A(start), .Z(n2892) );
  CNR2IXL U2147 ( .B(nst[2]), .A(n2892), .Z(N34) );
  CNIVXL U2148 ( .A(muordi), .Z(n2897) );
  CNR2XL U2149 ( .A(n2140), .B(n2895), .Z(n2167) );
  CNIVX1 U2150 ( .A(n922), .Z(n2894) );
  CNIVX1 U2151 ( .A(n2897), .Z(n2895) );
  CNIVX1 U2152 ( .A(n924), .Z(n2898) );
  CNIVX1 U2153 ( .A(n799), .Z(n2899) );
  CEOXL U2154 ( .A(opera2[27]), .B(opera2_63), .Z(n2807) );
  CNIVX1 U2155 ( .A(n800), .Z(n2900) );
  CENX1 U2156 ( .A(opera2[22]), .B(opera2_63), .Z(n2776) );
  CNIVX1 U2157 ( .A(n2776), .Z(n2901) );
  CEOXL U2158 ( .A(opera2[18]), .B(opera2_63), .Z(n2750) );
  CENX1 U2159 ( .A(opera2[16]), .B(opera2_63), .Z(n2738) );
  CNIVX1 U2160 ( .A(n2738), .Z(n2902) );
  CEOXL U2161 ( .A(n2737), .B(n2902), .Z(n2734) );
  CEOXL U2162 ( .A(opera2[15]), .B(opera2_63), .Z(n2731) );
  CENX1 U2163 ( .A(opera2[13]), .B(opera2_63), .Z(n2719) );
  CNIVX1 U2164 ( .A(n2719), .Z(n2903) );
  CNIVX1 U2165 ( .A(n813), .Z(n2904) );
  CEOXL U2166 ( .A(opera2[12]), .B(opera2_63), .Z(n2712) );
  CENX1 U2167 ( .A(opera2[10]), .B(opera2_63), .Z(n2700) );
  CNIVX1 U2168 ( .A(n2700), .Z(n2905) );
  CNIVX1 U2169 ( .A(n816), .Z(n2906) );
  CEOXL U2170 ( .A(opera2[9]), .B(opera2_63), .Z(n2693) );
  CENXL U2171 ( .A(opera2[7]), .B(opera2_63), .Z(n2681) );
  CEOXL U2172 ( .A(opera2[6]), .B(opera2_63), .Z(n2674) );
  CENX1 U2173 ( .A(opera2[4]), .B(opera2_63), .Z(n2662) );
  CNIVX1 U2174 ( .A(n2662), .Z(n2907) );
  CEOXL U2175 ( .A(opera2[3]), .B(opera2_63), .Z(n2655) );
  CENXL U2176 ( .A(opera2[1]), .B(opera2_63), .Z(n2642) );
  CNIVX1 U2177 ( .A(n825), .Z(n2908) );
  CNIVX1 U2178 ( .A(n806), .Z(n2909) );
  CENXL U2179 ( .A(opera2[19]), .B(opera2_63), .Z(n2757) );
  CNIVX1 U2180 ( .A(n801), .Z(n2910) );
  CEOXL U2181 ( .A(opera2[24]), .B(opera2_63), .Z(n2788) );
  CNIVX1 U2182 ( .A(n804), .Z(n2911) );
  CEOXL U2183 ( .A(opera2[21]), .B(opera2_63), .Z(n2769) );
  CNIVX1 U2184 ( .A(n856), .Z(n2912) );
  CENX1 U2185 ( .A(opera2[28]), .B(opera2_63), .Z(n2814) );
  CNIVX1 U2186 ( .A(n2814), .Z(n2913) );
  CNR3X1 U2187 ( .A(n2820), .B(n2814), .C(n2813), .Z(n2821) );
  COND1XL U2188 ( .A(n2998), .B(n3405), .C(n3404), .Z(n919) );
  CNR3X2 U2189 ( .A(n2643), .B(n2642), .C(n2649), .Z(n2650) );
  CNR2X1 U2190 ( .A(n2988), .B(n2936), .Z(n2927) );
  CANR1XL U2191 ( .A(n3427), .B(n3215), .C(n3214), .Z(n2929) );
  CENX1 U2192 ( .A(opera1[5]), .B(opera1[31]), .Z(n3137) );
  CNR2X1 U2193 ( .A(n3134), .B(n3139), .Z(n2931) );
  CANR11XL U2194 ( .A(n2867), .B(n3560), .C(n3532), .D(n3531), .Z(n3535) );
  CNR2IX1 U2195 ( .B(res_not_wire[42]), .A(n3443), .Z(n2956) );
  CND3XL U2196 ( .A(res_not_wire[44]), .B(n2956), .C(n3425), .Z(n3253) );
  CIVX2 U2197 ( .A(n3562), .Z(n3544) );
  CNR2X1 U2198 ( .A(n3416), .B(n2955), .Z(n2954) );
  CND2XL U2199 ( .A(n2933), .B(n3130), .Z(n3416) );
  COND2X1 U2200 ( .A(n3372), .B(n2033), .C(n3371), .D(n3370), .Z(n2934) );
  COND2XL U2201 ( .A(n3372), .B(n2033), .C(n3371), .D(n3370), .Z(n3540) );
  COND2XL U2202 ( .A(n3239), .B(n2113), .C(n3238), .D(n2929), .Z(n2935) );
  CNR3X2 U2203 ( .A(n2687), .B(n2681), .C(n2680), .Z(n2688) );
  CNR2X2 U2204 ( .A(n2661), .B(n2878), .Z(n2669) );
  CND2X1 U2205 ( .A(n2886), .B(res_not_wire[32]), .Z(n2936) );
  CNR3X1 U2206 ( .A(n2706), .B(n2700), .C(n2699), .Z(n2707) );
  CNR2X2 U2207 ( .A(n2737), .B(n2883), .Z(n2745) );
  CNR3X1 U2208 ( .A(n2725), .B(n2719), .C(n2718), .Z(n2726) );
  COND1XL U2209 ( .A(n3478), .B(n3476), .C(n2959), .Z(n3189) );
  CND2IX1 U2210 ( .B(n3296), .A(n3276), .Z(n3298) );
  COR2X1 U2211 ( .A(n3115), .B(n3138), .Z(n3134) );
  CANR4CXL U2212 ( .A(n2738), .B(n2737), .C(n2744), .D(n2745), .Z(n2741) );
  CENX1 U2213 ( .A(n3427), .B(n3426), .Z(n3428) );
  CND2X1 U2214 ( .A(n2669), .B(n2674), .Z(n2680) );
  CENX1 U2215 ( .A(opera1[7]), .B(opera1[31]), .Z(n3172) );
  CEOX1 U2216 ( .A(result[49]), .B(n3286), .Z(n3503) );
  CND3XL U2217 ( .A(n3565), .B(n3564), .C(n3563), .Z(n828) );
  CIVX2 U2218 ( .A(opera2[11]), .Z(n2943) );
  CEOXL U2219 ( .A(opera2[8]), .B(n2866), .Z(n2687) );
  CND3XL U2220 ( .A(n3442), .B(n3441), .C(n3440), .Z(n847) );
  CND3XL U2221 ( .A(n3500), .B(n3499), .C(n3498), .Z(n838) );
  CENX1 U2222 ( .A(opera1[11]), .B(n2877), .Z(n3201) );
  CENX1 U2223 ( .A(opera1[14]), .B(opera1[31]), .Z(n3234) );
  CEOXL U2224 ( .A(opera2[14]), .B(n2866), .Z(n2725) );
  CENX1 U2225 ( .A(opera1[15]), .B(opera1[31]), .Z(n3231) );
  CENX1 U2226 ( .A(opera1[17]), .B(opera1[31]), .Z(n3245) );
  CENX1 U2227 ( .A(opera1[23]), .B(opera1[31]), .Z(n3317) );
  CEOXL U2228 ( .A(opera2[5]), .B(n2866), .Z(n2668) );
  CND2IX2 U2229 ( .B(n2937), .A(c_inres), .Z(n3103) );
  CIVX2 U2230 ( .A(n3130), .Z(n2938) );
  CNR2X1 U2231 ( .A(n2995), .B(n2938), .Z(n2939) );
  CND2X1 U2232 ( .A(n2650), .B(n2655), .Z(n2661) );
  CANR4CXL U2233 ( .A(n2814), .B(n2813), .C(n2820), .D(n2821), .Z(n2817) );
  CND2XL U2234 ( .A(n2707), .B(n2712), .Z(n2718) );
  CND2XL U2235 ( .A(n2688), .B(n2693), .Z(n2699) );
  CENXL U2236 ( .A(n2826), .B(n2821), .Z(n2824) );
  CND2XL U2237 ( .A(n2764), .B(n2769), .Z(n2775) );
  CND2XL U2238 ( .A(n2783), .B(n2788), .Z(n2794) );
  CEOXL U2239 ( .A(n2813), .B(n2913), .Z(n2810) );
  CEOXL U2240 ( .A(n2794), .B(n2795), .Z(n2791) );
  CEOXL U2241 ( .A(n2775), .B(n2901), .Z(n2772) );
  CNR2XL U2242 ( .A(n3381), .B(n2029), .Z(n3382) );
  CNR2XL U2243 ( .A(n3335), .B(n2093), .Z(n3336) );
  CIVX1 U2244 ( .A(n3348), .Z(n3337) );
  CEOXL U2245 ( .A(n2769), .B(n2764), .Z(n2767) );
  CANR1XL U2246 ( .A(n3457), .B(n3466), .C(n3453), .Z(n3478) );
  CND2X1 U2247 ( .A(n3325), .B(n3324), .Z(n3326) );
  CEOXL U2248 ( .A(n2731), .B(n2726), .Z(n2729) );
  CND2XL U2249 ( .A(n2954), .B(n3196), .Z(n3433) );
  CEOXL U2250 ( .A(n3502), .B(n2940), .Z(n3506) );
  CAN2X1 U2251 ( .A(n3530), .B(n2949), .Z(n3531) );
  CANR4CXL U2252 ( .A(n2719), .B(n2718), .C(n2725), .D(n2726), .Z(n2722) );
  CEOXL U2253 ( .A(n2712), .B(n2707), .Z(n2710) );
  CIVX2 U2254 ( .A(n3558), .Z(n3530) );
  CANR4CXL U2255 ( .A(n2700), .B(n2699), .C(n2706), .D(n2707), .Z(n2703) );
  CNR3XL U2256 ( .A(n2250), .B(n2874), .C(n2137), .Z(n2259) );
  CANR4CXL U2257 ( .A(n2681), .B(n2680), .C(n2687), .D(n2688), .Z(n2684) );
  CEOXL U2258 ( .A(n3453), .B(n3458), .Z(n3459) );
  CND2X1 U2259 ( .A(n2745), .B(n2750), .Z(n2756) );
  CND2XL U2260 ( .A(n2815), .B(n2816), .Z(n796) );
  CND2IX1 U2261 ( .B(n2941), .A(n2823), .Z(n795) );
  CAOR2X2 U2262 ( .A(n3574), .B(result[31]), .C(result[30]), .D(n2871), .Z(
        n2941) );
  CND2XL U2263 ( .A(n2808), .B(n2809), .Z(n797) );
  CND2XL U2264 ( .A(n2796), .B(n2797), .Z(n799) );
  CND2XL U2265 ( .A(n2777), .B(n2778), .Z(n802) );
  CENX1 U2266 ( .A(n2943), .B(n2866), .Z(n2706) );
  CND2IX1 U2267 ( .B(n2944), .A(n2785), .Z(n801) );
  CAOR2X2 U2268 ( .A(n3574), .B(result[25]), .C(result[24]), .D(n2871), .Z(
        n2944) );
  COR2XL U2269 ( .A(n2961), .B(n3171), .Z(n3457) );
  COR2XL U2270 ( .A(n2964), .B(n3174), .Z(n3182) );
  COR2XL U2271 ( .A(n2957), .B(n3175), .Z(n3187) );
  CND2IX1 U2272 ( .B(n2945), .A(n2766), .Z(n804) );
  CAOR2X2 U2273 ( .A(n3574), .B(result[22]), .C(result[21]), .D(n2871), .Z(
        n2945) );
  CND2XL U2274 ( .A(n2751), .B(n2752), .Z(n806) );
  CENX1 U2275 ( .A(n2946), .B(n3386), .Z(n3545) );
  CND2XL U2276 ( .A(result[34]), .B(n2871), .Z(n2347) );
  COR2XL U2277 ( .A(n2962), .B(n3286), .Z(n3504) );
  COND3X1 U2278 ( .A(n3484), .B(n2870), .C(n3483), .D(n3482), .Z(n849) );
  COND3XL U2279 ( .A(n3435), .B(n3434), .C(n2867), .D(n3443), .Z(n3442) );
  COR2XL U2280 ( .A(n2963), .B(n3243), .Z(n3288) );
  CND2IXL U2281 ( .B(res_not_wire[42]), .A(n3443), .Z(n3444) );
  CNR2IXL U2282 ( .B(result[35]), .A(n3000), .Z(n3420) );
  CEOXL U2283 ( .A(n2661), .B(n2907), .Z(n2658) );
  CEOXL U2284 ( .A(n2699), .B(n2905), .Z(n2696) );
  CEOXL U2285 ( .A(n2642), .B(n2926), .Z(n2639) );
  CEOXL U2286 ( .A(n2680), .B(n2681), .Z(n2677) );
  CEOXL U2287 ( .A(n2693), .B(n2688), .Z(n2691) );
  CEOXL U2288 ( .A(n2718), .B(n2903), .Z(n2715) );
  CANR2XL U2289 ( .A(result[34]), .B(n3003), .C(n3002), .D(n2047), .Z(n2297)
         );
  CANR2XL U2290 ( .A(result[35]), .B(n3003), .C(n3002), .D(n2953), .Z(n2298)
         );
  CNR2IXL U2291 ( .B(result[33]), .A(n3001), .Z(n3126) );
  CMXI2XL U2292 ( .A0(n3002), .A1(n3003), .S(result[33]), .Z(n3568) );
  CMXI2XL U2293 ( .A0(n3002), .A1(n3003), .S(result[32]), .Z(n3570) );
  CIVXL U2294 ( .A(result[34]), .Z(n2047) );
  CIVXL U2295 ( .A(res_not_wire[6]), .Z(n2023) );
  CEOXL U2296 ( .A(n2750), .B(n2745), .Z(n2748) );
  CND2X1 U2297 ( .A(opera2[0]), .B(n2866), .Z(n2947) );
  CEOXL U2298 ( .A(c_inop2), .B(n2635), .Z(n2633) );
  CIVX2 U2299 ( .A(n3035), .Z(n3573) );
  CIVX2 U2300 ( .A(n2874), .Z(n3004) );
  CIVX2 U2301 ( .A(n2330), .Z(n3554) );
  CND2X1 U2302 ( .A(n2874), .B(n2247), .Z(n2178) );
  CND2X1 U2303 ( .A(n3586), .B(n2178), .Z(n2179) );
  COND1XL U2304 ( .A(n2149), .B(n2179), .C(n2178), .Z(n2187) );
  COND1XL U2305 ( .A(n2146), .B(n2179), .C(n2178), .Z(n2197) );
  COND1XL U2306 ( .A(n2150), .B(n2179), .C(n2178), .Z(n2177) );
  COND1XL U2307 ( .A(n2148), .B(n2179), .C(n2178), .Z(n2192) );
  COND1XL U2308 ( .A(n2144), .B(n2179), .C(n2178), .Z(n2209) );
  COND1XL U2309 ( .A(n2118), .B(n2179), .C(n2178), .Z(n2219) );
  COND1XL U2310 ( .A(n2130), .B(n2179), .C(n2178), .Z(n2214) );
  COND1XL U2311 ( .A(n2117), .B(n2179), .C(n2178), .Z(n2224) );
  COND1XL U2312 ( .A(n2105), .B(n2179), .C(n2178), .Z(n2229) );
  CNIVX1 U2313 ( .A(n2259), .Z(n3002) );
  CAN2X1 U2314 ( .A(n2247), .B(n2140), .Z(n2249) );
  CNR3XL U2315 ( .A(n2763), .B(n2757), .C(n2756), .Z(n2764) );
  CNR3XL U2316 ( .A(n2801), .B(n2795), .C(n2794), .Z(n2802) );
  CNR3XL U2317 ( .A(n2782), .B(n2776), .C(n2775), .Z(n2783) );
  CND2X1 U2318 ( .A(n3579), .B(n3574), .Z(n2330) );
  CANR1XL U2319 ( .A(n3134), .B(n3139), .C(n2931), .Z(n3135) );
  CENX1 U2320 ( .A(n2933), .B(n2116), .Z(n3117) );
  CNR2XL U2321 ( .A(n3373), .B(n2034), .Z(n3374) );
  CND2X1 U2322 ( .A(n2726), .B(n2731), .Z(n2737) );
  CNR2X1 U2323 ( .A(n3240), .B(n2040), .Z(n3241) );
  CNR2X1 U2324 ( .A(n3206), .B(n2044), .Z(n3207) );
  CEOXL U2325 ( .A(n3370), .B(n3371), .Z(n3342) );
  CNR2X1 U2326 ( .A(n3326), .B(n2035), .Z(n3327) );
  CNR2X1 U2327 ( .A(n3213), .B(n2115), .Z(n3214) );
  COND1XL U2328 ( .A(n2931), .B(n2882), .C(n3170), .Z(n3143) );
  CNR2X1 U2329 ( .A(n3137), .B(n3136), .Z(n3141) );
  CND2X1 U2330 ( .A(n3202), .B(n3203), .Z(n3437) );
  CENX1 U2331 ( .A(n2866), .B(n2003), .Z(n2826) );
  CND2X1 U2332 ( .A(n3378), .B(n3366), .Z(n3376) );
  CND2XL U2333 ( .A(n3369), .B(n3365), .Z(n3366) );
  CND2X1 U2334 ( .A(n3285), .B(n3284), .Z(n3300) );
  CND2X1 U2335 ( .A(n3298), .B(n3283), .Z(n3284) );
  CND2X1 U2336 ( .A(n3323), .B(n3282), .Z(n3321) );
  CND2XL U2337 ( .A(n3285), .B(n3281), .Z(n3282) );
  CND2XL U2338 ( .A(n3236), .B(n3231), .Z(n3232) );
  CNR2IX1 U2339 ( .B(n2779), .A(n3035), .Z(n3036) );
  CND2X1 U2340 ( .A(n3380), .B(n3379), .Z(n3381) );
  CND2XL U2341 ( .A(n3378), .B(n3377), .Z(n3379) );
  CND2XL U2342 ( .A(n3296), .B(n3295), .Z(n3297) );
  CND2XL U2343 ( .A(n3341), .B(n3334), .Z(n3335) );
  CND2XL U2344 ( .A(n3333), .B(n3332), .Z(n3334) );
  CND2XL U2345 ( .A(n3323), .B(n3322), .Z(n3324) );
  CND2XL U2346 ( .A(n3142), .B(n3105), .Z(n3115) );
  CNR2IXL U2347 ( .B(n2867), .A(n2954), .Z(n3147) );
  CNR2IXL U2348 ( .B(n2867), .A(n2956), .Z(n3445) );
  CND2XL U2349 ( .A(n3290), .B(n3247), .Z(n3286) );
  CND2XL U2350 ( .A(n3246), .B(n3245), .Z(n3247) );
  CND3XL U2351 ( .A(n3164), .B(n3163), .C(n3162), .Z(n856) );
  CND2X1 U2352 ( .A(n2252), .B(n3008), .Z(n3011) );
  CND2XL U2353 ( .A(n3106), .B(n3107), .Z(n3108) );
  CEOXL U2354 ( .A(n3529), .B(n3528), .Z(n2949) );
  CNR2IXL U2355 ( .B(n3153), .A(n3558), .Z(n3156) );
  CND3XL U2356 ( .A(n3129), .B(n3128), .C(n3127), .Z(n855) );
  CND2XL U2357 ( .A(n3530), .B(n3125), .Z(n3128) );
  CANR1XL U2358 ( .A(result[34]), .B(n3554), .C(n3126), .Z(n3127) );
  CND2XL U2359 ( .A(n3109), .B(n3108), .Z(n3154) );
  CNR2XL U2360 ( .A(n2950), .B(n3558), .Z(n3248) );
  CND2XL U2361 ( .A(n3454), .B(n3457), .Z(n3475) );
  CNR2IX1 U2362 ( .B(n3182), .A(n3475), .Z(n2951) );
  CEOXL U2363 ( .A(n3521), .B(n3522), .Z(n3523) );
  CEOXL U2364 ( .A(n3307), .B(n3308), .Z(n3309) );
  CNIVX1 U2365 ( .A(n2258), .Z(n3003) );
  CND2XL U2366 ( .A(n3287), .B(n3288), .Z(n3505) );
  CENX1 U2367 ( .A(n2935), .B(n3254), .Z(n3256) );
  CEOXL U2368 ( .A(n3494), .B(n3495), .Z(n3496) );
  CANR1XL U2369 ( .A(n2246), .B(n3005), .C(n2007), .Z(n2242) );
  CANR1XL U2370 ( .A(n2234), .B(n3005), .C(n2007), .Z(n2232) );
  CANR1XL U2371 ( .A(n2157), .B(n3005), .C(n2182), .Z(n2170) );
  CANR1XL U2372 ( .A(n2834), .B(n3576), .C(n2256), .Z(n3008) );
  CANR1XL U2373 ( .A(n2200), .B(n3005), .C(n2007), .Z(n2202) );
  CEOXL U2374 ( .A(n3485), .B(n3486), .Z(n3487) );
  COND2X1 U2375 ( .A(n2242), .B(n2120), .C(n2179), .D(n2243), .Z(n925) );
  CND2X1 U2376 ( .A(n3585), .B(n2120), .Z(n2243) );
  COND2X1 U2377 ( .A(n2232), .B(n2103), .C(n2179), .D(n2233), .Z(n929) );
  CEOX1 U2378 ( .A(n2756), .B(n2757), .Z(n2753) );
  CND2X1 U2379 ( .A(n2837), .B(n3586), .Z(n2247) );
  COND4CX1 U2380 ( .A(n2170), .B(n2171), .C(n2151), .D(n2172), .Z(n954) );
  CANR11XL U2381 ( .A(n2173), .B(n2151), .C(n3005), .D(n2008), .Z(n2172) );
  CND2XL U2382 ( .A(n3005), .B(n2156), .Z(n2171) );
  CEOXL U2383 ( .A(n2929), .B(n3238), .Z(n3219) );
  CEOXL U2384 ( .A(n3446), .B(n3447), .Z(n3448) );
  CENX1 U2385 ( .A(n2959), .B(n3479), .Z(n3480) );
  CANR1XL U2386 ( .A(n3478), .B(n3477), .C(n3476), .Z(n3479) );
  COND3XL U2387 ( .A(n3190), .B(n3189), .C(n3188), .D(n3187), .Z(n3191) );
  CND2X1 U2388 ( .A(n3584), .B(n2141), .Z(n2254) );
  CANR1XL U2389 ( .A(n2255), .B(n3586), .C(n2256), .Z(n2253) );
  CND2XL U2390 ( .A(n3454), .B(n3474), .Z(n3467) );
  CNIVXL U2391 ( .A(n3064), .Z(n2983) );
  CEOXL U2392 ( .A(n3079), .B(n2159), .Z(n3075) );
  CENX1 U2393 ( .A(n2982), .B(n3102), .Z(n3104) );
  CEOXL U2394 ( .A(n3088), .B(n2023), .Z(n3085) );
  CNR3XL U2395 ( .A(n3153), .B(n2250), .C(n3579), .Z(n3157) );
  CNIVXL U2396 ( .A(n3103), .Z(n2982) );
  CND4X1 U2397 ( .A(res_not_wire[40]), .B(n3196), .C(n2954), .D(n3434), .Z(
        n3443) );
  CEOX1 U2398 ( .A(result[39]), .B(n3174), .Z(n3453) );
  CEOX1 U2399 ( .A(result[43]), .B(n3209), .Z(n3446) );
  CEOX1 U2400 ( .A(result[42]), .B(n3206), .Z(n3436) );
  CNR2IXL U2401 ( .B(result[62]), .A(n3386), .Z(n3388) );
  CANR1XL U2402 ( .A(n3580), .B(n3386), .C(n3385), .Z(n3387) );
  CEOX1 U2403 ( .A(result[45]), .B(n3239), .Z(n3238) );
  CNR2IXL U2404 ( .B(n3406), .A(n3558), .Z(n3410) );
  CND2XL U2405 ( .A(n2330), .B(n3408), .Z(n3409) );
  CND2XL U2406 ( .A(n3574), .B(n3407), .Z(n3408) );
  CEOX1 U2407 ( .A(result[44]), .B(n3213), .Z(n3426) );
  CEOX1 U2408 ( .A(result[56]), .B(n3335), .Z(n3348) );
  CEOX1 U2409 ( .A(result[54]), .B(n3326), .Z(n3511) );
  CEOX1 U2410 ( .A(result[46]), .B(n3240), .Z(n3254) );
  CNR2IX1 U2411 ( .B(res_not_wire[40]), .A(n3433), .Z(n3435) );
  CND3XL U2412 ( .A(n3530), .B(n3203), .C(n3191), .Z(n3194) );
  CANR1XL U2413 ( .A(result[41]), .B(n3554), .C(n3192), .Z(n3193) );
  CANR1XL U2414 ( .A(n3425), .B(n2956), .C(res_not_wire[44]), .Z(n3224) );
  CND2XL U2415 ( .A(n3530), .B(n3219), .Z(n3222) );
  CND2XL U2416 ( .A(n3530), .B(n3301), .Z(n3304) );
  CANR1XL U2417 ( .A(result[53]), .B(n3554), .C(n3302), .Z(n3303) );
  CND2XL U2418 ( .A(n3530), .B(n3342), .Z(n3345) );
  CANR1XL U2419 ( .A(result[57]), .B(n3554), .C(n3343), .Z(n3344) );
  CANR1XL U2420 ( .A(result[60]), .B(n3554), .C(n3399), .Z(n3400) );
  CND2XL U2421 ( .A(n3530), .B(n3419), .Z(n3422) );
  CANR1XL U2422 ( .A(n3465), .B(n2954), .C(res_not_wire[38]), .Z(n3464) );
  CND2XL U2423 ( .A(n3530), .B(n3459), .Z(n3462) );
  CND2XL U2424 ( .A(n3530), .B(n3487), .Z(n3490) );
  CANR1XL U2425 ( .A(result[47]), .B(n3554), .C(n3488), .Z(n3489) );
  CANR1XL U2426 ( .A(result[45]), .B(n3554), .C(n3220), .Z(n3221) );
  CNR2IX1 U2427 ( .B(result[44]), .A(n3001), .Z(n3220) );
  CANR1XL U2428 ( .A(result[36]), .B(n3554), .C(n3420), .Z(n3421) );
  CANR1XL U2429 ( .A(result[39]), .B(n3554), .C(n3460), .Z(n3461) );
  CNR2IX1 U2430 ( .B(result[38]), .A(n3000), .Z(n3460) );
  CND2IX1 U2431 ( .B(n3558), .A(n3391), .Z(n3392) );
  CANR1XL U2432 ( .A(result[62]), .B(n3554), .C(n3548), .Z(n3549) );
  CENX1 U2433 ( .A(result[40]), .B(n3175), .Z(n2959) );
  COND3X1 U2434 ( .A(n3354), .B(n2868), .C(n3353), .D(n3352), .Z(n833) );
  CND2XL U2435 ( .A(n3530), .B(n3350), .Z(n3353) );
  CANR1XL U2436 ( .A(result[56]), .B(n3554), .C(n3351), .Z(n3352) );
  COND3XL U2437 ( .A(n2953), .B(n2330), .C(n2347), .D(n2348), .Z(n854) );
  COND3X1 U2438 ( .A(n3260), .B(n2870), .C(n3259), .D(n3258), .Z(n843) );
  CND2XL U2439 ( .A(n3530), .B(n3256), .Z(n3259) );
  CANR1XL U2440 ( .A(result[46]), .B(n3554), .C(n3257), .Z(n3258) );
  COND3X1 U2441 ( .A(n3313), .B(n2870), .C(n3312), .D(n3311), .Z(n837) );
  CND2XL U2442 ( .A(n3530), .B(n3309), .Z(n3312) );
  CANR1XL U2443 ( .A(result[52]), .B(n3554), .C(n3310), .Z(n3311) );
  COND3X1 U2444 ( .A(n3432), .B(n2998), .C(n3431), .D(n3430), .Z(n845) );
  CND2XL U2445 ( .A(n3530), .B(n3428), .Z(n3431) );
  CANR1XL U2446 ( .A(result[44]), .B(n3554), .C(n3429), .Z(n3430) );
  COND3X1 U2447 ( .A(n3472), .B(n2998), .C(n3471), .D(n3470), .Z(n851) );
  CND2XL U2448 ( .A(n3530), .B(n3468), .Z(n3471) );
  CANR1XL U2449 ( .A(result[38]), .B(n3554), .C(n3469), .Z(n3470) );
  CND2XL U2450 ( .A(n3530), .B(n3480), .Z(n3483) );
  CANR1XL U2451 ( .A(result[40]), .B(n3554), .C(n3481), .Z(n3482) );
  COND3X1 U2452 ( .A(n3510), .B(n2870), .C(n3509), .D(n3508), .Z(n839) );
  CND2XL U2453 ( .A(n3530), .B(n3506), .Z(n3509) );
  CANR1XL U2454 ( .A(result[50]), .B(n3554), .C(n3507), .Z(n3508) );
  CNR2XL U2455 ( .A(n3518), .B(n2960), .Z(n2992) );
  CANR2X1 U2456 ( .A(n2821), .B(n2003), .C(n2001), .D(n2866), .Z(n2833) );
  CNR2IX1 U2457 ( .B(result[61]), .A(n3000), .Z(n3548) );
  CNR2IX1 U2458 ( .B(result[36]), .A(n3001), .Z(n3148) );
  CNR2IX1 U2459 ( .B(result[40]), .A(n3001), .Z(n3192) );
  CNR2IX1 U2460 ( .B(result[48]), .A(n3001), .Z(n3250) );
  CNR2IX1 U2461 ( .B(result[45]), .A(n3001), .Z(n3257) );
  CNR2IX1 U2462 ( .B(result[47]), .A(n3001), .Z(n3268) );
  CNR2IX1 U2463 ( .B(result[52]), .A(n3000), .Z(n3302) );
  CNR2IX1 U2464 ( .B(result[51]), .A(n3000), .Z(n3310) );
  CNR2IX1 U2465 ( .B(result[56]), .A(n3001), .Z(n3343) );
  CNR2IX1 U2466 ( .B(result[55]), .A(n3000), .Z(n3351) );
  CNR2IX1 U2467 ( .B(result[59]), .A(n3000), .Z(n3399) );
  CNR2IX1 U2468 ( .B(result[43]), .A(n3000), .Z(n3429) );
  CNR2IX1 U2469 ( .B(result[41]), .A(n3000), .Z(n3439) );
  CNR2IX1 U2470 ( .B(result[42]), .A(n3000), .Z(n3449) );
  CNR2IX1 U2471 ( .B(result[37]), .A(n3001), .Z(n3469) );
  CNR2IX1 U2472 ( .B(result[39]), .A(n3000), .Z(n3481) );
  CNR2IX1 U2473 ( .B(result[46]), .A(n3001), .Z(n3488) );
  CNR2IX1 U2474 ( .B(result[50]), .A(n3001), .Z(n3497) );
  CNR2IX1 U2475 ( .B(result[49]), .A(n3000), .Z(n3507) );
  CNR2IX1 U2476 ( .B(result[53]), .A(n3001), .Z(n3514) );
  CNR2IX1 U2477 ( .B(result[54]), .A(n3000), .Z(n3524) );
  CNR2IX1 U2478 ( .B(result[57]), .A(n3000), .Z(n3541) );
  CND3XL U2479 ( .A(res_not_wire[38]), .B(n2954), .C(n3465), .Z(n3473) );
  CND3XL U2480 ( .A(n3517), .B(n3516), .C(n3515), .Z(n835) );
  CND2XL U2481 ( .A(n3530), .B(n3513), .Z(n3516) );
  CANR1XL U2482 ( .A(result[54]), .B(n3554), .C(n3514), .Z(n3515) );
  CANR1XL U2483 ( .A(result[58]), .B(n3554), .C(n3541), .Z(n3542) );
  CND2X1 U2484 ( .A(result[41]), .B(n3179), .Z(n3202) );
  CANR2XL U2485 ( .A(result[60]), .B(n2871), .C(result[61]), .D(n3554), .Z(
        n3565) );
  CND2XL U2486 ( .A(n3530), .B(n3523), .Z(n3526) );
  CANR1XL U2487 ( .A(result[55]), .B(n3554), .C(n3524), .Z(n3525) );
  CND3XL U2488 ( .A(n3271), .B(n3270), .C(n3269), .Z(n841) );
  CND2XL U2489 ( .A(n3530), .B(n3267), .Z(n3270) );
  CND2X1 U2490 ( .A(n3264), .B(n3263), .Z(n3271) );
  CANR1XL U2491 ( .A(result[48]), .B(n3554), .C(n3268), .Z(n3269) );
  CND2XL U2492 ( .A(n3530), .B(n3438), .Z(n3441) );
  CANR1XL U2493 ( .A(result[42]), .B(n3554), .C(n3439), .Z(n3440) );
  CND2X1 U2494 ( .A(n3445), .B(n3444), .Z(n3452) );
  CND2XL U2495 ( .A(n3530), .B(n3448), .Z(n3451) );
  CANR1XL U2496 ( .A(result[43]), .B(n3554), .C(n3449), .Z(n3450) );
  CND2XL U2497 ( .A(n3530), .B(n3496), .Z(n3499) );
  CND2X1 U2498 ( .A(n3493), .B(n3492), .Z(n3500) );
  CANR1XL U2499 ( .A(result[51]), .B(n3554), .C(n3497), .Z(n3498) );
  CANR1XL U2500 ( .A(result[59]), .B(n3554), .C(n3533), .Z(n3534) );
  CANR2XL U2501 ( .A(n3574), .B(result[15]), .C(result[14]), .D(n2871), .Z(
        n2720) );
  CNR2IX1 U2502 ( .B(result[62]), .A(n3000), .Z(n3357) );
  CENX1 U2503 ( .A(n134), .B(n2987), .Z(n3412) );
  CND2X1 U2504 ( .A(n3150), .B(n3149), .Z(n852) );
  CANR2XL U2505 ( .A(n3147), .B(n3146), .C(n3530), .D(n3145), .Z(n3150) );
  CANR1XL U2506 ( .A(result[37]), .B(n3554), .C(n3148), .Z(n3149) );
  CND2X1 U2507 ( .A(n3252), .B(n3251), .Z(n840) );
  CANR1XL U2508 ( .A(result[49]), .B(n3554), .C(n3250), .Z(n3251) );
  CND2X1 U2509 ( .A(n2630), .B(n2631), .Z(n825) );
  CANR2X1 U2510 ( .A(n3573), .B(n2633), .C(n2867), .D(n2634), .Z(n2631) );
  CANR2XL U2511 ( .A(n3574), .B(result[1]), .C(n2871), .D(result[0]), .Z(n2630) );
  CND2X1 U2512 ( .A(n2656), .B(n2657), .Z(n821) );
  CANR2X1 U2513 ( .A(n2658), .B(n3573), .C(n2867), .D(n3093), .Z(n2657) );
  CANR2XL U2514 ( .A(n3574), .B(result[5]), .C(result[4]), .D(n2871), .Z(n2656) );
  CANR2XL U2515 ( .A(n3574), .B(result[9]), .C(result[8]), .D(n2871), .Z(n2682) );
  CND2X1 U2516 ( .A(n2694), .B(n2695), .Z(n815) );
  CANR2X1 U2517 ( .A(n2696), .B(n3573), .C(n2869), .D(n3074), .Z(n2695) );
  CANR2XL U2518 ( .A(n3574), .B(result[11]), .C(result[10]), .D(n2871), .Z(
        n2694) );
  CND2X1 U2519 ( .A(n2708), .B(n2709), .Z(n813) );
  CANR2X1 U2520 ( .A(n2710), .B(n3573), .C(n2869), .D(n3067), .Z(n2709) );
  CANR2XL U2521 ( .A(n3574), .B(result[13]), .C(result[12]), .D(n2871), .Z(
        n2708) );
  CENX1 U2522 ( .A(n2147), .B(n3066), .Z(n3067) );
  CND2X1 U2523 ( .A(n2732), .B(n2733), .Z(n809) );
  CANR2X1 U2524 ( .A(n2734), .B(n3573), .C(n2867), .D(n3057), .Z(n2733) );
  CANR2XL U2525 ( .A(n3574), .B(result[17]), .C(result[16]), .D(n2871), .Z(
        n2732) );
  CENX1 U2526 ( .A(res_not_wire[16]), .B(n3056), .Z(n3057) );
  CND2X1 U2527 ( .A(n2746), .B(n2747), .Z(n807) );
  CANR2X1 U2528 ( .A(n2748), .B(n3573), .C(n2869), .D(n3049), .Z(n2747) );
  CANR2XL U2529 ( .A(n3574), .B(result[19]), .C(result[18]), .D(n2871), .Z(
        n2746) );
  CANR2XL U2530 ( .A(n3574), .B(result[21]), .C(result[20]), .D(n2871), .Z(
        n2758) );
  CND2X1 U2531 ( .A(n2770), .B(n2771), .Z(n803) );
  CANR2X1 U2532 ( .A(n2772), .B(n3573), .C(n2869), .D(n3039), .Z(n2771) );
  CANR2XL U2533 ( .A(n3574), .B(result[23]), .C(result[22]), .D(n2871), .Z(
        n2770) );
  CENX1 U2534 ( .A(n2952), .B(n2126), .Z(n3039) );
  CANR2X1 U2535 ( .A(n2786), .B(n3573), .C(n2869), .D(n3032), .Z(n2785) );
  CENX1 U2536 ( .A(n2124), .B(n3031), .Z(n3032) );
  CANR2XL U2537 ( .A(n3574), .B(result[27]), .C(result[26]), .D(n2871), .Z(
        n2796) );
  CANR2XL U2538 ( .A(n3574), .B(result[29]), .C(result[28]), .D(n2871), .Z(
        n2808) );
  CND2X1 U2539 ( .A(n2637), .B(n2638), .Z(n824) );
  CANR2X1 U2540 ( .A(n2639), .B(n3573), .C(n2869), .D(n3104), .Z(n2638) );
  CANR2XL U2541 ( .A(n3574), .B(result[2]), .C(result[1]), .D(n2871), .Z(n2637) );
  CND2X1 U2542 ( .A(n2651), .B(n2652), .Z(n822) );
  CANR2X1 U2543 ( .A(n2653), .B(n3573), .C(n2869), .D(n3095), .Z(n2652) );
  CANR2XL U2544 ( .A(n3574), .B(result[4]), .C(result[3]), .D(n2871), .Z(n2651) );
  CANR2XL U2545 ( .A(n3574), .B(result[6]), .C(result[5]), .D(n2871), .Z(n2663) );
  CND2X1 U2546 ( .A(n2675), .B(n2676), .Z(n818) );
  CANR2X1 U2547 ( .A(n2677), .B(n3573), .C(n2867), .D(n3084), .Z(n2676) );
  CANR2XL U2548 ( .A(n3574), .B(result[8]), .C(result[7]), .D(n2871), .Z(n2675) );
  CND2X1 U2549 ( .A(n2689), .B(n2690), .Z(n816) );
  CANR2X1 U2550 ( .A(n2691), .B(n3573), .C(n2867), .D(n3075), .Z(n2690) );
  CANR2XL U2551 ( .A(n3574), .B(result[10]), .C(result[9]), .D(n2871), .Z(
        n2689) );
  CANR2XL U2552 ( .A(n3574), .B(result[12]), .C(result[11]), .D(n2871), .Z(
        n2701) );
  CND2X1 U2553 ( .A(n2713), .B(n2714), .Z(n812) );
  CANR2X1 U2554 ( .A(n2715), .B(n3573), .C(n2869), .D(n3065), .Z(n2714) );
  CANR2XL U2555 ( .A(n3574), .B(result[14]), .C(result[13]), .D(n2871), .Z(
        n2713) );
  CND2X1 U2556 ( .A(n2727), .B(n2728), .Z(n810) );
  CANR2X1 U2557 ( .A(n2729), .B(n3573), .C(n2867), .D(n3059), .Z(n2728) );
  CANR2XL U2558 ( .A(n3574), .B(result[16]), .C(result[15]), .D(n2871), .Z(
        n2727) );
  CENX1 U2559 ( .A(n150), .B(n3058), .Z(n3059) );
  CANR2XL U2560 ( .A(n3574), .B(result[18]), .C(result[17]), .D(n2871), .Z(
        n2739) );
  CANR2X1 U2561 ( .A(n2753), .B(n3573), .C(n2869), .D(n3048), .Z(n2752) );
  CANR2XL U2562 ( .A(n3574), .B(result[20]), .C(result[19]), .D(n2871), .Z(
        n2751) );
  CENX1 U2563 ( .A(n146), .B(n2985), .Z(n3048) );
  CANR2XL U2564 ( .A(n3574), .B(result[24]), .C(result[23]), .D(n2871), .Z(
        n2777) );
  CND2X1 U2565 ( .A(n2789), .B(n2790), .Z(n800) );
  CANR2X1 U2566 ( .A(n2791), .B(n3573), .C(n2869), .D(n3030), .Z(n2790) );
  CANR2XL U2567 ( .A(n3574), .B(result[26]), .C(result[25]), .D(n2871), .Z(
        n2789) );
  CENX1 U2568 ( .A(n3029), .B(n3028), .Z(n3030) );
  CND2X1 U2569 ( .A(n2803), .B(n2804), .Z(n798) );
  CANR2XL U2570 ( .A(n3574), .B(result[28]), .C(result[27]), .D(n2871), .Z(
        n2803) );
  CENX1 U2571 ( .A(n138), .B(n3023), .Z(n3024) );
  CANR2XL U2572 ( .A(n3574), .B(result[30]), .C(result[29]), .D(n2871), .Z(
        n2815) );
  CND2X1 U2573 ( .A(n2670), .B(n2671), .Z(n819) );
  CANR2X1 U2574 ( .A(n2672), .B(n3573), .C(n2867), .D(n3085), .Z(n2671) );
  CANR2XL U2575 ( .A(n3574), .B(result[7]), .C(result[6]), .D(n2871), .Z(n2670) );
  CANR2XL U2576 ( .A(n3574), .B(result[3]), .C(result[2]), .D(n2871), .Z(n2644) );
  CND2X1 U2577 ( .A(n2151), .B(n2155), .Z(n2839) );
  COND1XL U2578 ( .A(n3004), .B(n2050), .C(n2838), .Z(n793) );
  COND1XL U2579 ( .A(n3004), .B(n2988), .C(n2293), .Z(n889) );
  CANR2X1 U2580 ( .A(result[30]), .B(n3003), .C(n3002), .D(n2068), .Z(n2293)
         );
  COND1XL U2581 ( .A(n3004), .B(n2090), .C(n2317), .Z(n865) );
  CANR2X1 U2582 ( .A(result[54]), .B(n3003), .C(n3002), .D(n2035), .Z(n2317)
         );
  CNR2IX1 U2583 ( .B(res_not_wire[38]), .A(n3004), .Z(n3273) );
  CNR2IX1 U2584 ( .B(res_not_wire[36]), .A(n3004), .Z(n3567) );
  CNR2IX1 U2585 ( .B(n2965), .A(n3004), .Z(n3569) );
  CNR2IX1 U2586 ( .B(res_not_wire[32]), .A(n3004), .Z(n3571) );
  CND3XL U2587 ( .A(n1119), .B(n2141), .C(n56), .Z(n2250) );
  COND1XL U2588 ( .A(i[12]), .B(n2179), .C(n2202), .Z(n2204) );
  CENX1 U2589 ( .A(opera1[18]), .B(n2877), .Z(n3289) );
  CENX1 U2590 ( .A(opera1[19]), .B(n2877), .Z(n3295) );
  CNR3XL U2591 ( .A(n3584), .B(n56), .C(n2141), .Z(n2834) );
  COND11XL U2592 ( .A(n2179), .B(i[12]), .C(n2200), .D(n2201), .Z(n942) );
  COND11X1 U2593 ( .A(n2179), .B(i[14]), .C(n2145), .D(n2205), .Z(n940) );
  COND4CX1 U2594 ( .A(n3005), .B(n2152), .C(n2204), .D(i[14]), .Z(n2205) );
  COND11X1 U2595 ( .A(n2179), .B(i[27]), .C(n2100), .D(n2237), .Z(n927) );
  CND2X1 U2596 ( .A(i[27]), .B(n2238), .Z(n2237) );
  COND11X1 U2597 ( .A(n2230), .B(n2106), .C(n2179), .D(n2231), .Z(n930) );
  COND4CX1 U2598 ( .A(n3005), .B(n2106), .C(n2229), .D(i[24]), .Z(n2231) );
  COND1XL U2599 ( .A(n164), .B(n3004), .C(n2264), .Z(n918) );
  CANR2X1 U2600 ( .A(result[1]), .B(n2258), .C(n3002), .D(n2067), .Z(n2264) );
  COND1XL U2601 ( .A(n3004), .B(n2159), .C(n2272), .Z(n910) );
  CANR2X1 U2602 ( .A(result[9]), .B(n3003), .C(n3002), .D(n2063), .Z(n2272) );
  COND1XL U2603 ( .A(n3004), .B(n2138), .C(n2257), .Z(n920) );
  CANR2X1 U2604 ( .A(result[0]), .B(n3003), .C(n3002), .D(n3579), .Z(n2257) );
  COND1XL U2605 ( .A(n150), .B(n3004), .C(n2278), .Z(n904) );
  CANR2X1 U2606 ( .A(result[15]), .B(n3003), .C(n3002), .D(n2060), .Z(n2278)
         );
  COND1XL U2607 ( .A(n160), .B(n3004), .C(n2268), .Z(n914) );
  CANR2X1 U2608 ( .A(result[5]), .B(n2258), .C(n2259), .D(n2065), .Z(n2268) );
  COND1XL U2609 ( .A(n3004), .B(n2133), .C(n2279), .Z(n903) );
  CANR2X1 U2610 ( .A(result[16]), .B(n3003), .C(n3002), .D(n2075), .Z(n2279)
         );
  COND1XL U2611 ( .A(n162), .B(n3004), .C(n2266), .Z(n916) );
  CANR2X1 U2612 ( .A(result[3]), .B(n3003), .C(n2259), .D(n2066), .Z(n2266) );
  COND1XL U2613 ( .A(n154), .B(n3004), .C(n2274), .Z(n908) );
  CANR2X1 U2614 ( .A(result[11]), .B(n3003), .C(n3002), .D(n2062), .Z(n2274)
         );
  COND1XL U2615 ( .A(n3004), .B(n3583), .C(n2283), .Z(n899) );
  CANR2X1 U2616 ( .A(result[20]), .B(n3003), .C(n3002), .D(n2073), .Z(n2283)
         );
  COND1XL U2617 ( .A(n3004), .B(n2126), .C(n2285), .Z(n897) );
  CANR2X1 U2618 ( .A(result[22]), .B(n3003), .C(n3002), .D(n2072), .Z(n2285)
         );
  COND1XL U2619 ( .A(n3004), .B(n2124), .C(n2287), .Z(n895) );
  CANR2X1 U2620 ( .A(result[24]), .B(n3003), .C(n3002), .D(n2071), .Z(n2287)
         );
  COND1XL U2621 ( .A(n148), .B(n3004), .C(n2280), .Z(n902) );
  CANR2X1 U2622 ( .A(result[17]), .B(n3003), .C(n3002), .D(n2059), .Z(n2280)
         );
  COND1XL U2623 ( .A(n3004), .B(n2116), .C(n2297), .Z(n885) );
  COND1XL U2624 ( .A(n3004), .B(n3582), .C(n2289), .Z(n893) );
  CANR2X1 U2625 ( .A(result[26]), .B(n3003), .C(n3002), .D(n2070), .Z(n2289)
         );
  COND1XL U2626 ( .A(n3004), .B(n2110), .C(n2291), .Z(n891) );
  CANR2X1 U2627 ( .A(result[28]), .B(n3003), .C(n3002), .D(n2069), .Z(n2291)
         );
  COND1XL U2628 ( .A(n138), .B(n3004), .C(n2290), .Z(n892) );
  CANR2X1 U2629 ( .A(result[27]), .B(n3003), .C(n3002), .D(n2054), .Z(n2290)
         );
  COND1XL U2630 ( .A(n136), .B(n3004), .C(n2292), .Z(n890) );
  CANR2X1 U2631 ( .A(result[29]), .B(n3003), .C(n3002), .D(n2053), .Z(n2292)
         );
  COND1XL U2632 ( .A(n126), .B(n3004), .C(n2302), .Z(n880) );
  CANR2X1 U2633 ( .A(result[39]), .B(n3003), .C(n3002), .D(n2964), .Z(n2302)
         );
  COND1XL U2634 ( .A(n3004), .B(n2096), .C(n2303), .Z(n879) );
  CANR2X1 U2635 ( .A(result[40]), .B(n3003), .C(n3002), .D(n2957), .Z(n2303)
         );
  COND1XL U2636 ( .A(n3004), .B(n2095), .C(n2305), .Z(n877) );
  CANR2X1 U2637 ( .A(result[42]), .B(n3003), .C(n3002), .D(n2044), .Z(n2305)
         );
  COND1XL U2638 ( .A(n3004), .B(n2094), .C(n2309), .Z(n873) );
  CANR2X1 U2639 ( .A(result[46]), .B(n3003), .C(n3002), .D(n2040), .Z(n2309)
         );
  COND1XL U2640 ( .A(n124), .B(n3004), .C(n2304), .Z(n878) );
  CANR2X1 U2641 ( .A(result[41]), .B(n3003), .C(n3002), .D(n2045), .Z(n2304)
         );
  COND1XL U2642 ( .A(n3004), .B(n2091), .C(n2315), .Z(n867) );
  CANR2X1 U2643 ( .A(result[52]), .B(n2258), .C(n3002), .D(n2098), .Z(n2315)
         );
  COND1XL U2644 ( .A(n3004), .B(n3581), .C(n2313), .Z(n869) );
  CANR2X1 U2645 ( .A(result[50]), .B(n3003), .C(n3002), .D(n2038), .Z(n2313)
         );
  COND1XL U2646 ( .A(n114), .B(n3004), .C(n2314), .Z(n868) );
  CANR2X1 U2647 ( .A(result[51]), .B(n2258), .C(n3002), .D(n2097), .Z(n2314)
         );
  COND1XL U2648 ( .A(n112), .B(n3004), .C(n2316), .Z(n866) );
  CANR2X1 U2649 ( .A(result[53]), .B(n3003), .C(n3002), .D(n2036), .Z(n2316)
         );
  COND1XL U2650 ( .A(n3004), .B(n2088), .C(n2311), .Z(n871) );
  CANR2X1 U2651 ( .A(result[48]), .B(n3003), .C(n3002), .D(n2963), .Z(n2311)
         );
  COND1XL U2652 ( .A(n3004), .B(n2085), .C(n2324), .Z(n858) );
  CANR2X1 U2653 ( .A(result[61]), .B(n2258), .C(n3002), .D(n2032), .Z(n2324)
         );
  COND1XL U2654 ( .A(n3004), .B(n3559), .C(n2323), .Z(n859) );
  CANR2X1 U2655 ( .A(result[60]), .B(n3003), .C(n3002), .D(n2029), .Z(n2323)
         );
  COND1XL U2656 ( .A(n106), .B(n3004), .C(n2322), .Z(n860) );
  CANR2X1 U2657 ( .A(result[59]), .B(n3003), .C(n3002), .D(n2086), .Z(n2322)
         );
  COND1XL U2658 ( .A(n146), .B(n3004), .C(n2282), .Z(n900) );
  CANR2X1 U2659 ( .A(result[19]), .B(n3003), .C(n2259), .D(n2058), .Z(n2282)
         );
  COND1XL U2660 ( .A(n142), .B(n3004), .C(n2286), .Z(n896) );
  CANR2X1 U2661 ( .A(result[23]), .B(n3003), .C(n3002), .D(n2056), .Z(n2286)
         );
  COND1XL U2662 ( .A(n144), .B(n3004), .C(n2284), .Z(n898) );
  CANR2X1 U2663 ( .A(result[21]), .B(n3003), .C(n2259), .D(n2057), .Z(n2284)
         );
  COND1XL U2664 ( .A(n130), .B(n3004), .C(n2298), .Z(n884) );
  COND1XL U2665 ( .A(n140), .B(n3004), .C(n2288), .Z(n894) );
  CANR2X1 U2666 ( .A(result[25]), .B(n3003), .C(n2259), .D(n2055), .Z(n2288)
         );
  COND1XL U2667 ( .A(n134), .B(n3004), .C(n2294), .Z(n888) );
  CANR2X1 U2668 ( .A(result[31]), .B(n3003), .C(n3002), .D(n2051), .Z(n2294)
         );
  COND1XL U2669 ( .A(n120), .B(n3004), .C(n2308), .Z(n874) );
  CANR2X1 U2670 ( .A(result[45]), .B(n3003), .C(n3002), .D(n2113), .Z(n2308)
         );
  COND1XL U2671 ( .A(n122), .B(n3004), .C(n2306), .Z(n876) );
  CANR2X1 U2672 ( .A(result[43]), .B(n2258), .C(n3002), .D(n2046), .Z(n2306)
         );
  COND1XL U2673 ( .A(n116), .B(n3004), .C(n2312), .Z(n870) );
  CANR2X1 U2674 ( .A(result[49]), .B(n3003), .C(n3002), .D(n2962), .Z(n2312)
         );
  COND1XL U2675 ( .A(n110), .B(n3004), .C(n2318), .Z(n864) );
  CANR2X1 U2676 ( .A(result[55]), .B(n3003), .C(n3002), .D(n2092), .Z(n2318)
         );
  COND1XL U2677 ( .A(n118), .B(n3004), .C(n2310), .Z(n872) );
  CANR2X1 U2678 ( .A(result[47]), .B(n2258), .C(n3002), .D(n2112), .Z(n2310)
         );
  COND1XL U2679 ( .A(n3004), .B(n2031), .C(n2325), .Z(n857) );
  CANR2X1 U2680 ( .A(result[62]), .B(n3003), .C(n3002), .D(n3580), .Z(n2325)
         );
  COND1XL U2681 ( .A(n3004), .B(n3536), .C(n2320), .Z(n862) );
  CANR2X1 U2682 ( .A(result[57]), .B(n3003), .C(n3002), .D(n2033), .Z(n2320)
         );
  COND1XL U2683 ( .A(n3004), .B(n3578), .C(n2321), .Z(n861) );
  CANR2X1 U2684 ( .A(result[58]), .B(n3003), .C(n3002), .D(n2034), .Z(n2321)
         );
  COND1XL U2685 ( .A(n128), .B(n3004), .C(n2300), .Z(n882) );
  CANR2X1 U2686 ( .A(result[37]), .B(n3003), .C(n3002), .D(n2042), .Z(n2300)
         );
  COND1XL U2687 ( .A(n3004), .B(n3577), .C(n2307), .Z(n875) );
  CANR2X1 U2688 ( .A(result[44]), .B(n3003), .C(n3002), .D(n2115), .Z(n2307)
         );
  COND1XL U2689 ( .A(n3004), .B(n3587), .C(n2319), .Z(n863) );
  CANR2X1 U2690 ( .A(result[56]), .B(n3003), .C(n3002), .D(n2093), .Z(n2319)
         );
  COND1XL U2691 ( .A(n158), .B(n3004), .C(n2270), .Z(n912) );
  CANR2X1 U2692 ( .A(result[7]), .B(n2258), .C(n3002), .D(n2064), .Z(n2270) );
  COND1XL U2693 ( .A(n3004), .B(n2023), .C(n2269), .Z(n913) );
  CANR2X1 U2694 ( .A(result[6]), .B(n3003), .C(n3002), .D(n2052), .Z(n2269) );
  COND1XL U2695 ( .A(n2170), .B(n2156), .C(n2183), .Z(n950) );
  CND4XL U2696 ( .A(i[1]), .B(n3005), .C(n2156), .D(i[0]), .Z(n2183) );
  COND1XL U2697 ( .A(n2005), .B(n2152), .C(n2203), .Z(n941) );
  COND1XL U2698 ( .A(n3004), .B(n2147), .C(n2275), .Z(n907) );
  CANR2X1 U2699 ( .A(result[12]), .B(n3003), .C(n3002), .D(n2077), .Z(n2275)
         );
  COND4CX1 U2700 ( .A(n2232), .B(n2235), .C(n2121), .D(n2236), .Z(n928) );
  CND2X1 U2701 ( .A(n3005), .B(n2103), .Z(n2235) );
  COND4CX1 U2702 ( .A(n2242), .B(n2244), .C(n2104), .D(n2245), .Z(n924) );
  CND2X1 U2703 ( .A(n3005), .B(n2120), .Z(n2244) );
  CND4X1 U2704 ( .A(i[29]), .B(n3005), .C(n2104), .D(n3585), .Z(n2245) );
  COND1XL U2705 ( .A(n3004), .B(n2125), .C(n2281), .Z(n901) );
  CANR2X1 U2706 ( .A(result[18]), .B(n3003), .C(n3002), .D(n2074), .Z(n2281)
         );
  CND3XL U2707 ( .A(n2175), .B(n2174), .C(n2176), .Z(n953) );
  COND4CX1 U2708 ( .A(n3005), .B(n2155), .C(n2177), .D(i[5]), .Z(n2176) );
  CND2X1 U2709 ( .A(valid), .B(n3575), .Z(n2252) );
  CNR2IX1 U2710 ( .B(n960), .A(n3004), .Z(n3118) );
  CANR2X1 U2711 ( .A(result[13]), .B(n3003), .C(n2259), .D(n2061), .Z(n2276)
         );
  CNR2IX1 U2712 ( .B(res_not_wire[10]), .A(n3004), .Z(n3119) );
  CANR2X1 U2713 ( .A(result[10]), .B(n3003), .C(n3002), .D(n2078), .Z(n2273)
         );
  CNR2IXL U2714 ( .B(res_not_wire[2]), .A(n3004), .Z(n3120) );
  CANR2X1 U2715 ( .A(result[2]), .B(n3003), .C(n2259), .D(n2081), .Z(n2265) );
  CNR2IX1 U2716 ( .B(res_not_wire[8]), .A(n3004), .Z(n3151) );
  CANR2X1 U2717 ( .A(result[8]), .B(n3003), .C(n3002), .D(n2079), .Z(n2271) );
  CNR2IX1 U2718 ( .B(res_not_wire[14]), .A(n3004), .Z(n3152) );
  CANR2X1 U2719 ( .A(result[14]), .B(n3003), .C(n2259), .D(n2076), .Z(n2277)
         );
  CNR2IX1 U2720 ( .B(res_not_wire[4]), .A(n3004), .Z(n3572) );
  CANR2X1 U2721 ( .A(result[4]), .B(n3003), .C(n3002), .D(n2080), .Z(n2267) );
  CND2X1 U2722 ( .A(n2188), .B(n2189), .Z(n947) );
  COND4CX1 U2723 ( .A(n3005), .B(n2163), .C(n2187), .D(i[7]), .Z(n2188) );
  CND2X1 U2724 ( .A(n2193), .B(n2194), .Z(n945) );
  COND4CX1 U2725 ( .A(n3005), .B(n2143), .C(n2192), .D(i[9]), .Z(n2193) );
  CND2X1 U2726 ( .A(n2198), .B(n2199), .Z(n943) );
  COND4CX1 U2727 ( .A(n3005), .B(n2154), .C(n2197), .D(i[11]), .Z(n2198) );
  CND2X1 U2728 ( .A(n2210), .B(n2211), .Z(n938) );
  COND4CX1 U2729 ( .A(n3005), .B(n2129), .C(n2209), .D(i[16]), .Z(n2210) );
  CND2X1 U2730 ( .A(n2220), .B(n2221), .Z(n934) );
  COND4CX1 U2731 ( .A(n3005), .B(n2123), .C(n2219), .D(i[20]), .Z(n2220) );
  CND2X1 U2732 ( .A(n2215), .B(n2216), .Z(n936) );
  COND4CX1 U2733 ( .A(n3005), .B(n2119), .C(n2214), .D(i[18]), .Z(n2215) );
  CND2X1 U2734 ( .A(n2225), .B(n2226), .Z(n932) );
  COND4CX1 U2735 ( .A(n3005), .B(n2122), .C(n2224), .D(i[22]), .Z(n2225) );
  CND2X1 U2736 ( .A(n2239), .B(n2240), .Z(n926) );
  COND4CX1 U2737 ( .A(n3005), .B(n2102), .C(n2238), .D(i[28]), .Z(n2239) );
  CENX1 U2738 ( .A(n960), .B(n2983), .Z(n3065) );
  CEOX1 U2739 ( .A(opera2[17]), .B(n2866), .Z(n2744) );
  CENX1 U2740 ( .A(opera1[20]), .B(n2877), .Z(n3283) );
  CENX1 U2741 ( .A(opera1[21]), .B(n2877), .Z(n3281) );
  CENX1 U2742 ( .A(opera1[22]), .B(n2877), .Z(n3322) );
  CENX1 U2743 ( .A(opera1[24]), .B(n2877), .Z(n3332) );
  COND1XL U2744 ( .A(i[0]), .B(n2179), .C(n2178), .Z(n2182) );
  COND11XL U2745 ( .A(n2179), .B(i[8]), .C(n2190), .D(n2191), .Z(n946) );
  CND2X1 U2746 ( .A(i[8]), .B(n2192), .Z(n2191) );
  COND11XL U2747 ( .A(n2179), .B(i[6]), .C(n2185), .D(n2186), .Z(n948) );
  CND2X1 U2748 ( .A(i[6]), .B(n2187), .Z(n2186) );
  CND2XL U2749 ( .A(i[1]), .B(n2182), .Z(n2181) );
  COND11XL U2750 ( .A(n2179), .B(i[4]), .C(n2180), .D(n2184), .Z(n949) );
  CND2X1 U2751 ( .A(i[4]), .B(n2177), .Z(n2184) );
  COND11XL U2752 ( .A(n2179), .B(i[10]), .C(n2195), .D(n2196), .Z(n944) );
  CND2X1 U2753 ( .A(i[10]), .B(n2197), .Z(n2196) );
  COND11XL U2754 ( .A(n2179), .B(i[15]), .C(n2207), .D(n2208), .Z(n939) );
  CND2X1 U2755 ( .A(i[15]), .B(n2209), .Z(n2208) );
  COND11XL U2756 ( .A(n2179), .B(i[19]), .C(n2217), .D(n2218), .Z(n935) );
  CND2X1 U2757 ( .A(i[19]), .B(n2219), .Z(n2218) );
  COND11XL U2758 ( .A(n2179), .B(i[21]), .C(n2222), .D(n2223), .Z(n933) );
  CND2X1 U2759 ( .A(i[21]), .B(n2224), .Z(n2223) );
  COND11XL U2760 ( .A(n2179), .B(i[17]), .C(n2212), .D(n2213), .Z(n937) );
  CND2X1 U2761 ( .A(i[17]), .B(n2214), .Z(n2213) );
  COND11XL U2762 ( .A(n2179), .B(i[23]), .C(n2227), .D(n2228), .Z(n931) );
  CND2X1 U2763 ( .A(i[23]), .B(n2229), .Z(n2228) );
  COND2XL U2764 ( .A(n2162), .B(n2178), .C(i[0]), .D(n2179), .Z(n952) );
  CND3XL U2765 ( .A(res_not_wire[38]), .B(n3465), .C(n3165), .Z(n3225) );
  CND3XL U2766 ( .A(n53), .B(n2178), .C(n56), .Z(n2174) );
  COND1XL U2767 ( .A(n2140), .B(n3576), .C(n2164), .Z(n957) );
  CANR2X1 U2768 ( .A(n3575), .B(n2016), .C(nst[0]), .D(n2166), .Z(n2164) );
  COND1XL U2769 ( .A(n2250), .B(n2101), .C(n2251), .Z(n921) );
  CANR2X1 U2770 ( .A(n3575), .B(n2016), .C(nst[2]), .D(n2166), .Z(n2251) );
  CIVX2 U2771 ( .A(result[61]), .Z(n2032) );
  CENX1 U2772 ( .A(n3014), .B(res_not_wire[10]), .Z(n3074) );
  CENX1 U2773 ( .A(opera1[25]), .B(n2877), .Z(n3340) );
  CENX1 U2774 ( .A(opera1[26]), .B(n2877), .Z(n3367) );
  CENX1 U2775 ( .A(opera1[27]), .B(n2877), .Z(n3365) );
  CENX1 U2776 ( .A(opera1[28]), .B(n2877), .Z(n3377) );
  CENX1 U2777 ( .A(opera1[29]), .B(n2877), .Z(n3364) );
  CEOX1 U2778 ( .A(opera2[20]), .B(n2866), .Z(n2763) );
  CEOX1 U2779 ( .A(opera2[23]), .B(n2866), .Z(n2782) );
  COND1XL U2780 ( .A(n2016), .B(n2049), .C(n2249), .Z(n922) );
  CIVX2 U2781 ( .A(result[62]), .Z(n3580) );
  CENX1 U2782 ( .A(n162), .B(n3094), .Z(n3095) );
  CENX1 U2783 ( .A(n158), .B(n3083), .Z(n3084) );
  CENX1 U2784 ( .A(opera1[30]), .B(n2877), .Z(n3385) );
  CEOX1 U2785 ( .A(opera2[26]), .B(n2866), .Z(n2801) );
  CEOX1 U2786 ( .A(n2866), .B(n2877), .Z(n3121) );
  CNR2X1 U2787 ( .A(n2892), .B(nst[0]), .Z(n55) );
  CND2X1 U2788 ( .A(result[63]), .B(n2871), .Z(n3404) );
  CANR1XL U2789 ( .A(result[63]), .B(n3554), .C(n3357), .Z(n3393) );
  CANR2X1 U2790 ( .A(result[63]), .B(n3003), .C(n3002), .D(n3588), .Z(n2838)
         );
  CIVXL U2791 ( .A(n2241), .Z(n2100) );
  COND1XL U2792 ( .A(n2241), .B(n2179), .C(n2178), .Z(n2238) );
  CENX1 U2793 ( .A(opera1[4]), .B(opera1[31]), .Z(n3139) );
  CND2X1 U2794 ( .A(n3535), .B(n3534), .Z(n830) );
  CNR3XL U2795 ( .A(n3501), .B(n116), .C(n3581), .Z(n2979) );
  CIVX2 U2796 ( .A(n3103), .Z(n2980) );
  CND2X1 U2797 ( .A(n2720), .B(n2721), .Z(n811) );
  CIVX2 U2798 ( .A(n3064), .Z(n2981) );
  CANR2X1 U2799 ( .A(n2767), .B(n3573), .C(n2869), .D(n3041), .Z(n2766) );
  COND2X1 U2800 ( .A(n3239), .B(n2113), .C(n3238), .D(n3237), .Z(n3255) );
  CNR2X1 U2801 ( .A(n3139), .B(n3138), .Z(n3140) );
  CNR2IXL U2802 ( .B(res_not_wire[18]), .A(n3052), .Z(n2985) );
  CNR2XL U2803 ( .A(n3018), .B(n2988), .Z(n2987) );
  CEOXL U2804 ( .A(n2674), .B(n2669), .Z(n2672) );
  CEOXL U2805 ( .A(n2655), .B(n2650), .Z(n2653) );
  CEOXL U2806 ( .A(n2788), .B(n2783), .Z(n2786) );
  CEOXL U2807 ( .A(n2807), .B(n2802), .Z(n2805) );
  CANR4CXL U2808 ( .A(n2795), .B(n2794), .C(n2801), .D(n2802), .Z(n2798) );
  CANR4CXL U2809 ( .A(n2776), .B(n2775), .C(n2782), .D(n2783), .Z(n2779) );
  CANR4CXL U2810 ( .A(n2662), .B(n2661), .C(n2668), .D(n2669), .Z(n2665) );
  CANR4CXL U2811 ( .A(n2642), .B(n2926), .C(n2649), .D(n2650), .Z(n2646) );
  CIVX2 U2812 ( .A(n3518), .Z(n2989) );
  CND2X1 U2813 ( .A(n3520), .B(n3519), .Z(n3527) );
  CNR2IXL U2814 ( .B(res_not_wire[52]), .A(n3314), .Z(n2990) );
  CND2IX2 U2815 ( .B(n112), .A(n2997), .Z(n3518) );
  CANR4CXL U2816 ( .A(n2757), .B(n2756), .C(n2763), .D(n2764), .Z(n2760) );
  CEOXL U2817 ( .A(n3556), .B(n3555), .Z(n3557) );
  CNR2IXL U2818 ( .B(n2951), .A(n3186), .Z(n3190) );
  CENX1 U2819 ( .A(opera1[3]), .B(opera1[31]), .Z(n3138) );
  CENX1 U2820 ( .A(opera1[2]), .B(opera1[31]), .Z(n3136) );
  CENX1 U2821 ( .A(result[63]), .B(n3390), .Z(n3391) );
  COND1XL U2822 ( .A(n3417), .B(n3180), .C(n3181), .Z(n3455) );
  CND2XL U2823 ( .A(result[36]), .B(n2846), .Z(n3181) );
  CND2X1 U2824 ( .A(res_not_wire[14]), .B(n960), .Z(n2996) );
  CENX1 U2825 ( .A(n3403), .B(n2050), .Z(n3405) );
  CND3XL U2826 ( .A(n3562), .B(n3561), .C(n2867), .Z(n3563) );
  CND3XL U2827 ( .A(n2869), .B(n3538), .C(n3537), .Z(n3543) );
  COND1XL U2828 ( .A(n2984), .B(n3587), .C(n3536), .Z(n3537) );
  CNR2IXL U2829 ( .B(n3033), .A(n2998), .Z(n3038) );
  COND1XL U2830 ( .A(n3077), .B(n158), .C(n3076), .Z(n3078) );
  COND1XL U2831 ( .A(n2982), .B(n164), .C(n3096), .Z(n3097) );
  CND2IXL U2832 ( .B(res_not_wire[58]), .A(n3538), .Z(n3532) );
  CND2IXL U2833 ( .B(res_not_wire[48]), .A(n3226), .Z(n3249) );
  CNR2IXL U2834 ( .B(n3025), .A(n2868), .Z(n3027) );
  CANR1XL U2835 ( .A(n1053), .B(n3544), .C(res_not_wire[62]), .Z(n3395) );
  COND3XL U2836 ( .A(n2990), .B(n2888), .C(n2869), .D(n3518), .Z(n3517) );
  CANR11XL U2837 ( .A(n3063), .B(n3062), .C(n2867), .D(n2881), .Z(n2721) );
  CND3XL U2838 ( .A(n2869), .B(n3098), .C(n3097), .Z(n3101) );
  CNR2IXL U2839 ( .B(n3018), .A(n2870), .Z(n3020) );
  CNR3XL U2840 ( .A(n2874), .B(n1061), .C(n2250), .Z(n2258) );
  CND2IXL U2841 ( .B(n2868), .A(n3416), .Z(n3423) );
  CNR2IXL U2842 ( .B(n2867), .A(n3261), .Z(n3264) );
  COND3X1 U2843 ( .A(n3402), .B(n2868), .C(n3401), .D(n3400), .Z(n829) );
  CND3XL U2844 ( .A(n2867), .B(n3070), .C(n3069), .Z(n3073) );
  CND3XL U2845 ( .A(n2867), .B(n3088), .C(n3087), .Z(n3091) );
  CND2IXL U2846 ( .B(n146), .A(n2985), .Z(n3042) );
  CNR2IXL U2847 ( .B(n2867), .A(n2992), .Z(n3520) );
  CNR2IXL U2848 ( .B(n2867), .A(n2979), .Z(n3493) );
  CANR1XL U2849 ( .A(res_not_wire[34]), .B(n2933), .C(n3415), .Z(n3424) );
  CANR11XL U2850 ( .A(n2867), .B(n3501), .C(n3249), .D(n3248), .Z(n3252) );
  CANR11XL U2851 ( .A(n2869), .B(n3161), .C(n3160), .D(n3159), .Z(n3162) );
  COND1XL U2852 ( .A(n3501), .B(n116), .C(n3581), .Z(n3492) );
  CND3XL U2853 ( .A(n2867), .B(n3052), .C(n3051), .Z(n3055) );
  COND1XL U2854 ( .A(n3560), .B(n106), .C(n3559), .Z(n3561) );
  CND3XL U2855 ( .A(n2869), .B(n3079), .C(n3078), .Z(n3082) );
  CND3XL U2856 ( .A(n2869), .B(n3044), .C(n3043), .Z(n3047) );
  COND1XL U2857 ( .A(n2983), .B(n3061), .C(n3060), .Z(n3062) );
  CND2IXL U2858 ( .B(n134), .A(n2987), .Z(n3158) );
  CNR2XL U2859 ( .A(n2987), .B(n2998), .Z(n3017) );
  COND1XL U2860 ( .A(n3029), .B(n140), .C(n3582), .Z(n3026) );
  CIVXL U2861 ( .A(n2179), .Z(n3005) );
  CAN2X1 U2862 ( .A(n53), .B(n56), .Z(n3006) );
  CND2IX1 U2863 ( .B(n1119), .A(n3006), .Z(n3015) );
  CIVX2 U2864 ( .A(n3015), .Z(n3575) );
  CIVX2 U2865 ( .A(n2895), .Z(n3576) );
  CIVX2 U2866 ( .A(n2250), .Z(n3586) );
  CIVX2 U2867 ( .A(n3009), .Z(n2169) );
  CIVX2 U2868 ( .A(result[63]), .Z(n3588) );
  CIVX2 U2869 ( .A(n1056), .Z(n2050) );
  CND2IX1 U2870 ( .B(n2247), .A(n3009), .Z(n3010) );
  CND2IX1 U2871 ( .B(n2250), .A(n3553), .Z(n3012) );
  CIVX2 U2872 ( .A(n3012), .Z(n3574) );
  CIVX2 U2873 ( .A(n140), .Z(n3028) );
  CIVX2 U2874 ( .A(res_not_wire[26]), .Z(n3582) );
  CIVX2 U2875 ( .A(n144), .Z(n3040) );
  CIVX2 U2876 ( .A(n164), .Z(n3102) );
  CIVX2 U2877 ( .A(n3098), .Z(n3094) );
  CIVX2 U2878 ( .A(n3079), .Z(n3013) );
  CND2X2 U2879 ( .A(res_not_wire[12]), .B(n3066), .Z(n3064) );
  CANR2X1 U2880 ( .A(n2824), .B(n3573), .C(n3017), .D(n3016), .Z(n2823) );
  CANR2X1 U2881 ( .A(n2817), .B(n3573), .C(n3020), .D(n3019), .Z(n2816) );
  CANR2X1 U2882 ( .A(n2810), .B(n3573), .C(n2867), .D(n3022), .Z(n2809) );
  CANR2X1 U2883 ( .A(n2805), .B(n3573), .C(n2867), .D(n3024), .Z(n2804) );
  CANR2X1 U2884 ( .A(n2798), .B(n3573), .C(n3027), .D(n3026), .Z(n2797) );
  CIVX2 U2885 ( .A(res_not_wire[22]), .Z(n2126) );
  CND2IX1 U2886 ( .B(res_not_wire[20]), .A(n3042), .Z(n3043) );
  CIVX2 U2887 ( .A(n2760), .Z(n3045) );
  CND2IX1 U2888 ( .B(n3045), .A(n3573), .Z(n3046) );
  CIVX2 U2889 ( .A(n2741), .Z(n3053) );
  CND2IX1 U2890 ( .B(n3053), .A(n3573), .Z(n3054) );
  CIVX2 U2891 ( .A(n960), .Z(n3061) );
  CIVX2 U2892 ( .A(res_not_wire[14]), .Z(n3060) );
  CIVX2 U2893 ( .A(n2703), .Z(n3071) );
  CND2IX1 U2894 ( .B(n3071), .A(n3573), .Z(n3072) );
  CIVX2 U2895 ( .A(res_not_wire[8]), .Z(n3076) );
  CIVX2 U2896 ( .A(n2684), .Z(n3080) );
  CND2IX1 U2897 ( .B(n3080), .A(n3573), .Z(n3081) );
  CIVX2 U2898 ( .A(n2665), .Z(n3089) );
  CND2IX1 U2899 ( .B(n3089), .A(n3573), .Z(n3090) );
  CIVX2 U2900 ( .A(res_not_wire[2]), .Z(n3096) );
  CIVX2 U2901 ( .A(n2646), .Z(n3099) );
  CND2IX1 U2902 ( .B(n3099), .A(n3573), .Z(n3100) );
  CIVX2 U2903 ( .A(res_not_wire[34]), .Z(n2116) );
  CENX1 U2904 ( .A(opera1[31]), .B(opera1[1]), .Z(n3106) );
  CIVX2 U2905 ( .A(n3136), .Z(n3105) );
  CIVX2 U2906 ( .A(n3112), .Z(n3124) );
  CIVX2 U2907 ( .A(n3407), .Z(n3406) );
  CIVX2 U2908 ( .A(n3153), .Z(n3111) );
  CIVX2 U2909 ( .A(n3123), .Z(n3114) );
  CND2IX1 U2910 ( .B(result[34]), .A(n3112), .Z(n3113) );
  COND4CX1 U2911 ( .A(result[34]), .B(n3124), .C(n3114), .D(n3113), .Z(n3132)
         );
  CANR2X1 U2912 ( .A(n2867), .B(n3117), .C(n3530), .D(n3116), .Z(n2348) );
  CIVX2 U2913 ( .A(n1053), .Z(n2085) );
  CIVX2 U2914 ( .A(result[60]), .Z(n2029) );
  CIVX2 U2915 ( .A(result[59]), .Z(n2086) );
  CIVX2 U2916 ( .A(result[58]), .Z(n2034) );
  CIVX2 U2917 ( .A(res_not_wire[58]), .Z(n3578) );
  CIVX2 U2918 ( .A(result[57]), .Z(n2033) );
  CIVX2 U2919 ( .A(result[56]), .Z(n2093) );
  CIVX2 U2920 ( .A(res_not_wire[56]), .Z(n3587) );
  CIVX2 U2921 ( .A(result[55]), .Z(n2092) );
  CIVX2 U2922 ( .A(result[54]), .Z(n2035) );
  CIVX2 U2923 ( .A(result[53]), .Z(n2036) );
  CIVX2 U2924 ( .A(result[52]), .Z(n2098) );
  CIVX2 U2925 ( .A(res_not_wire[52]), .Z(n2091) );
  CIVX2 U2926 ( .A(result[51]), .Z(n2097) );
  CIVX2 U2927 ( .A(result[50]), .Z(n2038) );
  CIVX2 U2928 ( .A(res_not_wire[50]), .Z(n3581) );
  CIVX2 U2929 ( .A(result[47]), .Z(n2112) );
  CIVX2 U2930 ( .A(result[46]), .Z(n2040) );
  CIVX2 U2931 ( .A(res_not_wire[46]), .Z(n2094) );
  CIVX2 U2932 ( .A(result[45]), .Z(n2113) );
  CIVX2 U2933 ( .A(result[44]), .Z(n2115) );
  CIVX2 U2934 ( .A(res_not_wire[44]), .Z(n3577) );
  CIVX2 U2935 ( .A(result[43]), .Z(n2046) );
  CIVX2 U2936 ( .A(result[42]), .Z(n2044) );
  CIVX2 U2937 ( .A(res_not_wire[40]), .Z(n2096) );
  CIVX2 U2938 ( .A(res_not_wire[28]), .Z(n2110) );
  CIVX2 U2939 ( .A(res_not_wire[20]), .Z(n3583) );
  CIVX2 U2940 ( .A(res_not_wire[16]), .Z(n2133) );
  CIVX2 U2941 ( .A(n2246), .Z(n3585) );
  CND2IX1 U2942 ( .B(n3118), .A(n2276), .Z(n906) );
  CND2IX1 U2943 ( .B(n3119), .A(n2273), .Z(n909) );
  CND2IX1 U2944 ( .B(n3120), .A(n2265), .Z(n917) );
  CEO3X1 U2945 ( .A(n2047), .B(n3124), .C(n3123), .Z(n3125) );
  CIVX2 U2946 ( .A(n130), .Z(n3415) );
  CND2IX1 U2947 ( .B(result[37]), .A(n3143), .Z(n3144) );
  CENX1 U2948 ( .A(n3455), .B(n3456), .Z(n3145) );
  CND2IX1 U2949 ( .B(n3151), .A(n2271), .Z(n911) );
  CND2IX1 U2950 ( .B(n3152), .A(n2277), .Z(n905) );
  CND2IX1 U2951 ( .B(n2928), .A(n3554), .Z(n3164) );
  CENX1 U2952 ( .A(result[33]), .B(n3154), .Z(n3155) );
  CMXI2X1 U2953 ( .A0(n3157), .A1(n3156), .S(n3155), .Z(n3163) );
  CND2IX1 U2954 ( .B(res_not_wire[32]), .A(n3158), .Z(n3160) );
  CIVX2 U2955 ( .A(n128), .Z(n3465) );
  CENX1 U2956 ( .A(n3433), .B(n2096), .Z(n3195) );
  CIVX2 U2957 ( .A(n3170), .Z(n3167) );
  CIVX2 U2958 ( .A(n3182), .Z(n3476) );
  CIVX2 U2959 ( .A(n3178), .Z(n3177) );
  CIVX2 U2960 ( .A(n3180), .Z(n3418) );
  CIVX2 U2961 ( .A(n3186), .Z(n3183) );
  CND2X1 U2962 ( .A(n3185), .B(n3184), .Z(n3203) );
  COND3X1 U2963 ( .A(n3195), .B(n2868), .C(n3194), .D(n3193), .Z(n848) );
  CIVX2 U2964 ( .A(n122), .Z(n3425) );
  CIVX2 U2965 ( .A(n3225), .Z(n3196) );
  CIVX2 U2966 ( .A(n124), .Z(n3434) );
  CND2IX1 U2967 ( .B(n2868), .A(n3253), .Z(n3223) );
  CIVX2 U2968 ( .A(n3204), .Z(n3198) );
  CIVX2 U2969 ( .A(n3205), .Z(n3200) );
  CIVX2 U2970 ( .A(n3201), .Z(n3199) );
  CIVX2 U2971 ( .A(n3436), .Z(n3208) );
  CIVX2 U2972 ( .A(n3426), .Z(n3215) );
  CIVX2 U2973 ( .A(n3218), .Z(n3217) );
  COND3X1 U2974 ( .A(n3224), .B(n3223), .C(n3222), .D(n3221), .Z(n844) );
  CIVX2 U2975 ( .A(n3226), .Z(n3261) );
  CND2X2 U2976 ( .A(res_not_wire[48]), .B(n3261), .Z(n3501) );
  CIVX2 U2977 ( .A(n3234), .Z(n3227) );
  CIVX2 U2978 ( .A(n3231), .Z(n3228) );
  CIVX2 U2979 ( .A(n3233), .Z(n3230) );
  CIVX2 U2980 ( .A(n3254), .Z(n3242) );
  CIVX2 U2981 ( .A(n3245), .Z(n3244) );
  CENX1 U2982 ( .A(n120), .B(n3253), .Z(n3260) );
  CMXI2X1 U2983 ( .A0(n3002), .A1(n2258), .S(result[38]), .Z(n3272) );
  CND2IX1 U2984 ( .B(n3273), .A(n3272), .Z(n881) );
  CIVX2 U2985 ( .A(n114), .Z(n3306) );
  CIVX2 U2986 ( .A(n3290), .Z(n3275) );
  CIVX2 U2987 ( .A(n3289), .Z(n3274) );
  CIVX2 U2988 ( .A(n3295), .Z(n3276) );
  CIVX2 U2989 ( .A(n3298), .Z(n3278) );
  CIVX2 U2990 ( .A(n3283), .Z(n3277) );
  CIVX2 U2991 ( .A(n3285), .Z(n3280) );
  CIVX2 U2992 ( .A(n3281), .Z(n3279) );
  CIVX2 U2993 ( .A(n3291), .Z(n3292) );
  COND3X1 U2994 ( .A(n3305), .B(n2868), .C(n3304), .D(n3303), .Z(n836) );
  CIVX2 U2995 ( .A(n110), .Z(n3347) );
  CIVX2 U2996 ( .A(n3323), .Z(n3316) );
  CIVX2 U2997 ( .A(n3322), .Z(n3315) );
  CIVX2 U2998 ( .A(n3318), .Z(n3319) );
  CIVX2 U2999 ( .A(n3511), .Z(n3328) );
  COND2X2 U3000 ( .A(n3329), .B(n2092), .C(n3522), .D(n3521), .Z(n3349) );
  CIVX2 U3001 ( .A(n3333), .Z(n3331) );
  CIVX2 U3002 ( .A(n3332), .Z(n3330) );
  CIVX2 U3003 ( .A(n3341), .Z(n3339) );
  CIVX2 U3004 ( .A(n3340), .Z(n3338) );
  COND3X1 U3005 ( .A(n3346), .B(n2870), .C(n3345), .D(n3344), .Z(n832) );
  CIVX2 U3006 ( .A(res_not_wire[60]), .Z(n3559) );
  CIVX2 U3007 ( .A(n3538), .Z(n3355) );
  CAN2X1 U3008 ( .A(res_not_wire[62]), .B(n1053), .Z(n3356) );
  CND2X2 U3009 ( .A(n3544), .B(n3356), .Z(n3403) );
  CIVX2 U3010 ( .A(n3368), .Z(n3359) );
  CIVX2 U3011 ( .A(n3367), .Z(n3358) );
  CIVX2 U3012 ( .A(n3369), .Z(n3361) );
  CIVX2 U3013 ( .A(n3365), .Z(n3360) );
  CIVX2 U3014 ( .A(n3378), .Z(n3363) );
  CIVX2 U3015 ( .A(n3377), .Z(n3362) );
  CIVX2 U3016 ( .A(n3545), .Z(n3389) );
  CIVX2 U3017 ( .A(n3539), .Z(n3375) );
  CIVX2 U3018 ( .A(n3396), .Z(n3383) );
  COND2X2 U3019 ( .A(n3384), .B(n2032), .C(n3555), .D(n3556), .Z(n3546) );
  CND2IX1 U3020 ( .B(n3558), .A(n3398), .Z(n3401) );
  CANR2X1 U3021 ( .A(n2829), .B(n3573), .C(n2869), .D(n3412), .Z(n3413) );
  CENX1 U3022 ( .A(n3418), .B(n3417), .Z(n3419) );
  COND3X1 U3023 ( .A(n3424), .B(n3423), .C(n3422), .D(n3421), .Z(n853) );
  CENX1 U3024 ( .A(n2956), .B(n3425), .Z(n3432) );
  CENX1 U3025 ( .A(n3437), .B(n3436), .Z(n3438) );
  CND2IX1 U3026 ( .B(n3456), .A(n3455), .Z(n3474) );
  COND3X1 U3027 ( .A(n3464), .B(n3463), .C(n3462), .D(n3461), .Z(n850) );
  CENX1 U3028 ( .A(n3467), .B(n3466), .Z(n3468) );
  CENX1 U3029 ( .A(n126), .B(n3473), .Z(n3484) );
  CND2IX1 U3030 ( .B(n3475), .A(n3474), .Z(n3477) );
  COND3X1 U3031 ( .A(n3491), .B(n2998), .C(n3490), .D(n3489), .Z(n842) );
  CIVX2 U3032 ( .A(n1093), .Z(n3536) );
  CENX1 U3033 ( .A(n3546), .B(n3545), .Z(n3547) );
  COND3X1 U3034 ( .A(n3552), .B(n2998), .C(n3550), .D(n3549), .Z(n827) );
  CND2IX1 U3035 ( .B(n3558), .A(n3557), .Z(n3564) );
  CMXI2X1 U3036 ( .A0(n2259), .A1(n2258), .S(result[36]), .Z(n3566) );
  CND2IX1 U3037 ( .B(n3567), .A(n3566), .Z(n883) );
  CND2IX1 U3038 ( .B(n3569), .A(n3568), .Z(n886) );
  CND2IX1 U3039 ( .B(n3571), .A(n3570), .Z(n887) );
  CND2IX1 U3040 ( .B(n3572), .A(n2267), .Z(n915) );
endmodule

